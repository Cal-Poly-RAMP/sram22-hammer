*SPICE NETLIST
* OPEN SOURCE CONVERSION PRELUDE (SPECTRE)

.SUBCKT sky130_fd_pr__special_nfet_pass d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b npass l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__special_nfet_latch d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b npd l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__nfet_01v8 d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b nshort l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__pfet_01v8 d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b pshort l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__special_pfet_pass d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b ppu l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__pfet_01v8_hvt d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b phighvt l='l' w='w' mult='mult'
.ENDS

.SUBCKT sky130_fd_pr__nfet_01v8_lvt d g s b
.PARAM w=1.0 l=1.0 mult=1
M0 d g s b nlowvt l='l' w='w' mult='mult'
.ENDS
* circuit.Package sramgen_sramgen_sram_32x32m8w32_replica_v1
* Written by SpiceNetlister
* 

.SUBCKT hierarchical_decoder_nand_1 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_inv_2 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder 
+ vdd gnd addr[1] addr[0] addr_b[1] addr_b[0] decode[3] decode[2] decode[1] decode[0] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_3 
+ gnd vdd addr_b[1] addr_b[0] decode_b[0] 
+ hierarchical_decoder_nand_1 
* No parameters

xinv_4 
+ gnd vdd decode_b[0] decode[0] 
+ hierarchical_decoder_inv_2 
* No parameters

xnand_5 
+ gnd vdd addr_b[1] addr[0] decode_b[1] 
+ hierarchical_decoder_nand_1 
* No parameters

xinv_6 
+ gnd vdd decode_b[1] decode[1] 
+ hierarchical_decoder_inv_2 
* No parameters

xnand_7 
+ gnd vdd addr[1] addr_b[0] decode_b[2] 
+ hierarchical_decoder_nand_1 
* No parameters

xinv_8 
+ gnd vdd decode_b[2] decode[2] 
+ hierarchical_decoder_inv_2 
* No parameters

xnand_9 
+ gnd vdd addr[1] addr[0] decode_b[3] 
+ hierarchical_decoder_nand_1 
* No parameters

xinv_10 
+ gnd vdd decode_b[3] decode[3] 
+ hierarchical_decoder_inv_2 
* No parameters

.ENDS

.SUBCKT column_decoder_nand_1 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder_inv_2 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder 
+ vdd gnd addr[2] addr[1] addr[0] addr_b[2] addr_b[1] addr_b[0] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_3 
+ gnd vdd addr_b[2] addr_b[1] addr_b[0] decode_b[0] 
+ column_decoder_nand_1 
* No parameters

xinv_4 
+ gnd vdd decode_b[0] decode[0] 
+ column_decoder_inv_2 
* No parameters

xnand_5 
+ gnd vdd addr_b[2] addr_b[1] addr[0] decode_b[1] 
+ column_decoder_nand_1 
* No parameters

xinv_6 
+ gnd vdd decode_b[1] decode[1] 
+ column_decoder_inv_2 
* No parameters

xnand_7 
+ gnd vdd addr_b[2] addr[1] addr_b[0] decode_b[2] 
+ column_decoder_nand_1 
* No parameters

xinv_8 
+ gnd vdd decode_b[2] decode[2] 
+ column_decoder_inv_2 
* No parameters

xnand_9 
+ gnd vdd addr_b[2] addr[1] addr[0] decode_b[3] 
+ column_decoder_nand_1 
* No parameters

xinv_10 
+ gnd vdd decode_b[3] decode[3] 
+ column_decoder_inv_2 
* No parameters

xnand_11 
+ gnd vdd addr[2] addr_b[1] addr_b[0] decode_b[4] 
+ column_decoder_nand_1 
* No parameters

xinv_12 
+ gnd vdd decode_b[4] decode[4] 
+ column_decoder_inv_2 
* No parameters

xnand_13 
+ gnd vdd addr[2] addr_b[1] addr[0] decode_b[5] 
+ column_decoder_nand_1 
* No parameters

xinv_14 
+ gnd vdd decode_b[5] decode[5] 
+ column_decoder_inv_2 
* No parameters

xnand_15 
+ gnd vdd addr[2] addr[1] addr_b[0] decode_b[6] 
+ column_decoder_nand_1 
* No parameters

xinv_16 
+ gnd vdd decode_b[6] decode[6] 
+ column_decoder_inv_2 
* No parameters

xnand_17 
+ gnd vdd addr[2] addr[1] addr[0] decode_b[7] 
+ column_decoder_nand_1 
* No parameters

xinv_18 
+ gnd vdd decode_b[7] decode[7] 
+ column_decoder_inv_2 
* No parameters

.ENDS

.SUBCKT wordline_driver_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ wordline_driver_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ wordline_driver_and2_inv 
* No parameters

.ENDS

.SUBCKT wordline_driver 
+ vdd vss din wl_en wl 

xand2 
+ din wl_en wl vdd vss 
+ wordline_driver_and2 
* No parameters

.ENDS

.SUBCKT wordline_driver_array 
+ vdd vss din[3] din[2] din[1] din[0] wl_en wl[3] wl[2] wl[1] wl[0] 

xwl_driver_0 
+ vdd vss din[0] wl_en wl[0] 
+ wordline_driver 
* No parameters

xwl_driver_1 
+ vdd vss din[1] wl_en wl[1] 
+ wordline_driver 
* No parameters

xwl_driver_2 
+ vdd vss din[2] wl_en wl[2] 
+ wordline_driver 
* No parameters

xwl_driver_3 
+ vdd vss din[3] wl_en wl[3] 
+ wordline_driver 
* No parameters

.ENDS

.SUBCKT bitcell_array 
+ vdd vss bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[3] wl[2] wl[1] wl[0] vnb vpb rbl rbr 

xbitcell_0_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_0 
+ vdd vdd vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_1 
+ rbl rbr vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_2 
+ bl[0] br[0] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_3 
+ bl[1] br[1] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_4 
+ bl[2] br[2] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_5 
+ bl[3] br[3] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_6 
+ bl[4] br[4] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_7 
+ bl[5] br[5] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_8 
+ bl[6] br[6] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_9 
+ bl[7] br[7] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_10 
+ bl[8] br[8] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_11 
+ bl[9] br[9] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_12 
+ bl[10] br[10] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_13 
+ bl[11] br[11] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_14 
+ bl[12] br[12] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_15 
+ bl[13] br[13] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_16 
+ bl[14] br[14] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_17 
+ bl[15] br[15] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_18 
+ bl[16] br[16] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_19 
+ bl[17] br[17] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_20 
+ bl[18] br[18] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_21 
+ bl[19] br[19] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_22 
+ bl[20] br[20] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_23 
+ bl[21] br[21] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_24 
+ bl[22] br[22] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_25 
+ bl[23] br[23] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_26 
+ bl[24] br[24] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_27 
+ bl[25] br[25] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_28 
+ bl[26] br[26] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_29 
+ bl[27] br[27] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_30 
+ bl[28] br[28] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_31 
+ bl[29] br[29] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_32 
+ bl[30] br[30] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_33 
+ bl[31] br[31] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_34 
+ bl[32] br[32] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_35 
+ bl[33] br[33] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_36 
+ bl[34] br[34] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_37 
+ bl[35] br[35] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_38 
+ bl[36] br[36] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_39 
+ bl[37] br[37] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_40 
+ bl[38] br[38] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_41 
+ bl[39] br[39] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_42 
+ bl[40] br[40] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_43 
+ bl[41] br[41] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_44 
+ bl[42] br[42] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_45 
+ bl[43] br[43] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_46 
+ bl[44] br[44] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_47 
+ bl[45] br[45] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_48 
+ bl[46] br[46] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_49 
+ bl[47] br[47] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_50 
+ bl[48] br[48] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_51 
+ bl[49] br[49] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_52 
+ bl[50] br[50] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_53 
+ bl[51] br[51] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_54 
+ bl[52] br[52] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_55 
+ bl[53] br[53] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_56 
+ bl[54] br[54] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_57 
+ bl[55] br[55] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_58 
+ bl[56] br[56] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_59 
+ bl[57] br[57] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_60 
+ bl[58] br[58] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_61 
+ bl[59] br[59] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_62 
+ bl[60] br[60] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_63 
+ bl[61] br[61] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_64 
+ bl[62] br[62] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_65 
+ bl[63] br[63] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_66 
+ bl[64] br[64] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_67 
+ bl[65] br[65] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_68 
+ bl[66] br[66] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_69 
+ bl[67] br[67] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_70 
+ bl[68] br[68] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_71 
+ bl[69] br[69] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_72 
+ bl[70] br[70] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_73 
+ bl[71] br[71] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_74 
+ bl[72] br[72] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_75 
+ bl[73] br[73] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_76 
+ bl[74] br[74] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_77 
+ bl[75] br[75] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_78 
+ bl[76] br[76] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_79 
+ bl[77] br[77] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_80 
+ bl[78] br[78] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_81 
+ bl[79] br[79] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_82 
+ bl[80] br[80] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_83 
+ bl[81] br[81] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_84 
+ bl[82] br[82] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_85 
+ bl[83] br[83] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_86 
+ bl[84] br[84] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_87 
+ bl[85] br[85] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_88 
+ bl[86] br[86] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_89 
+ bl[87] br[87] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_90 
+ bl[88] br[88] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_91 
+ bl[89] br[89] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_92 
+ bl[90] br[90] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_93 
+ bl[91] br[91] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_94 
+ bl[92] br[92] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_95 
+ bl[93] br[93] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_96 
+ bl[94] br[94] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_97 
+ bl[95] br[95] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_98 
+ bl[96] br[96] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_99 
+ bl[97] br[97] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_100 
+ bl[98] br[98] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_101 
+ bl[99] br[99] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_102 
+ bl[100] br[100] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_103 
+ bl[101] br[101] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_104 
+ bl[102] br[102] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_105 
+ bl[103] br[103] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_106 
+ bl[104] br[104] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_107 
+ bl[105] br[105] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_108 
+ bl[106] br[106] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_109 
+ bl[107] br[107] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_110 
+ bl[108] br[108] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_111 
+ bl[109] br[109] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_112 
+ bl[110] br[110] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_113 
+ bl[111] br[111] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_114 
+ bl[112] br[112] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_115 
+ bl[113] br[113] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_116 
+ bl[114] br[114] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_117 
+ bl[115] br[115] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_118 
+ bl[116] br[116] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_119 
+ bl[117] br[117] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_120 
+ bl[118] br[118] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_121 
+ bl[119] br[119] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_122 
+ bl[120] br[120] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_123 
+ bl[121] br[121] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_124 
+ bl[122] br[122] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_125 
+ bl[123] br[123] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_126 
+ bl[124] br[124] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_127 
+ bl[125] br[125] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_128 
+ bl[126] br[126] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_129 
+ bl[127] br[127] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_130 
+ bl[128] br[128] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_131 
+ bl[129] br[129] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_132 
+ bl[130] br[130] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_133 
+ bl[131] br[131] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_134 
+ bl[132] br[132] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_135 
+ bl[133] br[133] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_136 
+ bl[134] br[134] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_137 
+ bl[135] br[135] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_138 
+ bl[136] br[136] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_139 
+ bl[137] br[137] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_140 
+ bl[138] br[138] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_141 
+ bl[139] br[139] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_142 
+ bl[140] br[140] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_143 
+ bl[141] br[141] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_144 
+ bl[142] br[142] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_145 
+ bl[143] br[143] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_146 
+ bl[144] br[144] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_147 
+ bl[145] br[145] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_148 
+ bl[146] br[146] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_149 
+ bl[147] br[147] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_150 
+ bl[148] br[148] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_151 
+ bl[149] br[149] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_152 
+ bl[150] br[150] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_153 
+ bl[151] br[151] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_154 
+ bl[152] br[152] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_155 
+ bl[153] br[153] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_156 
+ bl[154] br[154] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_157 
+ bl[155] br[155] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_158 
+ bl[156] br[156] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_159 
+ bl[157] br[157] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_160 
+ bl[158] br[158] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_161 
+ bl[159] br[159] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_162 
+ bl[160] br[160] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_163 
+ bl[161] br[161] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_164 
+ bl[162] br[162] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_165 
+ bl[163] br[163] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_166 
+ bl[164] br[164] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_167 
+ bl[165] br[165] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_168 
+ bl[166] br[166] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_169 
+ bl[167] br[167] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_170 
+ bl[168] br[168] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_171 
+ bl[169] br[169] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_172 
+ bl[170] br[170] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_173 
+ bl[171] br[171] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_174 
+ bl[172] br[172] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_175 
+ bl[173] br[173] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_176 
+ bl[174] br[174] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_177 
+ bl[175] br[175] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_178 
+ bl[176] br[176] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_179 
+ bl[177] br[177] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_180 
+ bl[178] br[178] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_181 
+ bl[179] br[179] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_182 
+ bl[180] br[180] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_183 
+ bl[181] br[181] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_184 
+ bl[182] br[182] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_185 
+ bl[183] br[183] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_186 
+ bl[184] br[184] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_187 
+ bl[185] br[185] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_188 
+ bl[186] br[186] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_189 
+ bl[187] br[187] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_190 
+ bl[188] br[188] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_191 
+ bl[189] br[189] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_192 
+ bl[190] br[190] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_193 
+ bl[191] br[191] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_194 
+ bl[192] br[192] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_195 
+ bl[193] br[193] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_196 
+ bl[194] br[194] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_197 
+ bl[195] br[195] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_198 
+ bl[196] br[196] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_199 
+ bl[197] br[197] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_200 
+ bl[198] br[198] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_201 
+ bl[199] br[199] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_202 
+ bl[200] br[200] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_203 
+ bl[201] br[201] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_204 
+ bl[202] br[202] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_205 
+ bl[203] br[203] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_206 
+ bl[204] br[204] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_207 
+ bl[205] br[205] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_208 
+ bl[206] br[206] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_209 
+ bl[207] br[207] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_210 
+ bl[208] br[208] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_211 
+ bl[209] br[209] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_212 
+ bl[210] br[210] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_213 
+ bl[211] br[211] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_214 
+ bl[212] br[212] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_215 
+ bl[213] br[213] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_216 
+ bl[214] br[214] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_217 
+ bl[215] br[215] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_218 
+ bl[216] br[216] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_219 
+ bl[217] br[217] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_220 
+ bl[218] br[218] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_221 
+ bl[219] br[219] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_222 
+ bl[220] br[220] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_223 
+ bl[221] br[221] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_224 
+ bl[222] br[222] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_225 
+ bl[223] br[223] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_226 
+ bl[224] br[224] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_227 
+ bl[225] br[225] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_228 
+ bl[226] br[226] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_229 
+ bl[227] br[227] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_230 
+ bl[228] br[228] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_231 
+ bl[229] br[229] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_232 
+ bl[230] br[230] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_233 
+ bl[231] br[231] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_234 
+ bl[232] br[232] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_235 
+ bl[233] br[233] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_236 
+ bl[234] br[234] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_237 
+ bl[235] br[235] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_238 
+ bl[236] br[236] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_239 
+ bl[237] br[237] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_240 
+ bl[238] br[238] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_241 
+ bl[239] br[239] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_242 
+ bl[240] br[240] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_243 
+ bl[241] br[241] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_244 
+ bl[242] br[242] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_245 
+ bl[243] br[243] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_246 
+ bl[244] br[244] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_247 
+ bl[245] br[245] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_248 
+ bl[246] br[246] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_249 
+ bl[247] br[247] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_250 
+ bl[248] br[248] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_251 
+ bl[249] br[249] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_252 
+ bl[250] br[250] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_253 
+ bl[251] br[251] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_254 
+ bl[252] br[252] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_255 
+ bl[253] br[253] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_256 
+ bl[254] br[254] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_257 
+ bl[255] br[255] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_258 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_259 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_0 
+ vdd vdd vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_1 
+ rbl rbr vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_2 
+ bl[0] br[0] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_3 
+ bl[1] br[1] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_4 
+ bl[2] br[2] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_5 
+ bl[3] br[3] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_6 
+ bl[4] br[4] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_7 
+ bl[5] br[5] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_8 
+ bl[6] br[6] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_9 
+ bl[7] br[7] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_10 
+ bl[8] br[8] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_11 
+ bl[9] br[9] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_12 
+ bl[10] br[10] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_13 
+ bl[11] br[11] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_14 
+ bl[12] br[12] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_15 
+ bl[13] br[13] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_16 
+ bl[14] br[14] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_17 
+ bl[15] br[15] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_18 
+ bl[16] br[16] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_19 
+ bl[17] br[17] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_20 
+ bl[18] br[18] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_21 
+ bl[19] br[19] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_22 
+ bl[20] br[20] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_23 
+ bl[21] br[21] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_24 
+ bl[22] br[22] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_25 
+ bl[23] br[23] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_26 
+ bl[24] br[24] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_27 
+ bl[25] br[25] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_28 
+ bl[26] br[26] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_29 
+ bl[27] br[27] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_30 
+ bl[28] br[28] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_31 
+ bl[29] br[29] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_32 
+ bl[30] br[30] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_33 
+ bl[31] br[31] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_34 
+ bl[32] br[32] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_35 
+ bl[33] br[33] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_36 
+ bl[34] br[34] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_37 
+ bl[35] br[35] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_38 
+ bl[36] br[36] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_39 
+ bl[37] br[37] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_40 
+ bl[38] br[38] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_41 
+ bl[39] br[39] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_42 
+ bl[40] br[40] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_43 
+ bl[41] br[41] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_44 
+ bl[42] br[42] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_45 
+ bl[43] br[43] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_46 
+ bl[44] br[44] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_47 
+ bl[45] br[45] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_48 
+ bl[46] br[46] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_49 
+ bl[47] br[47] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_50 
+ bl[48] br[48] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_51 
+ bl[49] br[49] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_52 
+ bl[50] br[50] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_53 
+ bl[51] br[51] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_54 
+ bl[52] br[52] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_55 
+ bl[53] br[53] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_56 
+ bl[54] br[54] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_57 
+ bl[55] br[55] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_58 
+ bl[56] br[56] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_59 
+ bl[57] br[57] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_60 
+ bl[58] br[58] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_61 
+ bl[59] br[59] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_62 
+ bl[60] br[60] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_63 
+ bl[61] br[61] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_64 
+ bl[62] br[62] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_65 
+ bl[63] br[63] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_66 
+ bl[64] br[64] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_67 
+ bl[65] br[65] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_68 
+ bl[66] br[66] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_69 
+ bl[67] br[67] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_70 
+ bl[68] br[68] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_71 
+ bl[69] br[69] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_72 
+ bl[70] br[70] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_73 
+ bl[71] br[71] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_74 
+ bl[72] br[72] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_75 
+ bl[73] br[73] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_76 
+ bl[74] br[74] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_77 
+ bl[75] br[75] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_78 
+ bl[76] br[76] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_79 
+ bl[77] br[77] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_80 
+ bl[78] br[78] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_81 
+ bl[79] br[79] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_82 
+ bl[80] br[80] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_83 
+ bl[81] br[81] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_84 
+ bl[82] br[82] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_85 
+ bl[83] br[83] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_86 
+ bl[84] br[84] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_87 
+ bl[85] br[85] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_88 
+ bl[86] br[86] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_89 
+ bl[87] br[87] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_90 
+ bl[88] br[88] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_91 
+ bl[89] br[89] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_92 
+ bl[90] br[90] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_93 
+ bl[91] br[91] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_94 
+ bl[92] br[92] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_95 
+ bl[93] br[93] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_96 
+ bl[94] br[94] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_97 
+ bl[95] br[95] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_98 
+ bl[96] br[96] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_99 
+ bl[97] br[97] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_100 
+ bl[98] br[98] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_101 
+ bl[99] br[99] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_102 
+ bl[100] br[100] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_103 
+ bl[101] br[101] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_104 
+ bl[102] br[102] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_105 
+ bl[103] br[103] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_106 
+ bl[104] br[104] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_107 
+ bl[105] br[105] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_108 
+ bl[106] br[106] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_109 
+ bl[107] br[107] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_110 
+ bl[108] br[108] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_111 
+ bl[109] br[109] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_112 
+ bl[110] br[110] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_113 
+ bl[111] br[111] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_114 
+ bl[112] br[112] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_115 
+ bl[113] br[113] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_116 
+ bl[114] br[114] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_117 
+ bl[115] br[115] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_118 
+ bl[116] br[116] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_119 
+ bl[117] br[117] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_120 
+ bl[118] br[118] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_121 
+ bl[119] br[119] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_122 
+ bl[120] br[120] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_123 
+ bl[121] br[121] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_124 
+ bl[122] br[122] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_125 
+ bl[123] br[123] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_126 
+ bl[124] br[124] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_127 
+ bl[125] br[125] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_128 
+ bl[126] br[126] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_129 
+ bl[127] br[127] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_130 
+ bl[128] br[128] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_131 
+ bl[129] br[129] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_132 
+ bl[130] br[130] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_133 
+ bl[131] br[131] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_134 
+ bl[132] br[132] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_135 
+ bl[133] br[133] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_136 
+ bl[134] br[134] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_137 
+ bl[135] br[135] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_138 
+ bl[136] br[136] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_139 
+ bl[137] br[137] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_140 
+ bl[138] br[138] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_141 
+ bl[139] br[139] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_142 
+ bl[140] br[140] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_143 
+ bl[141] br[141] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_144 
+ bl[142] br[142] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_145 
+ bl[143] br[143] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_146 
+ bl[144] br[144] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_147 
+ bl[145] br[145] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_148 
+ bl[146] br[146] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_149 
+ bl[147] br[147] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_150 
+ bl[148] br[148] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_151 
+ bl[149] br[149] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_152 
+ bl[150] br[150] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_153 
+ bl[151] br[151] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_154 
+ bl[152] br[152] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_155 
+ bl[153] br[153] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_156 
+ bl[154] br[154] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_157 
+ bl[155] br[155] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_158 
+ bl[156] br[156] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_159 
+ bl[157] br[157] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_160 
+ bl[158] br[158] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_161 
+ bl[159] br[159] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_162 
+ bl[160] br[160] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_163 
+ bl[161] br[161] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_164 
+ bl[162] br[162] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_165 
+ bl[163] br[163] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_166 
+ bl[164] br[164] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_167 
+ bl[165] br[165] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_168 
+ bl[166] br[166] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_169 
+ bl[167] br[167] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_170 
+ bl[168] br[168] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_171 
+ bl[169] br[169] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_172 
+ bl[170] br[170] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_173 
+ bl[171] br[171] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_174 
+ bl[172] br[172] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_175 
+ bl[173] br[173] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_176 
+ bl[174] br[174] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_177 
+ bl[175] br[175] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_178 
+ bl[176] br[176] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_179 
+ bl[177] br[177] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_180 
+ bl[178] br[178] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_181 
+ bl[179] br[179] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_182 
+ bl[180] br[180] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_183 
+ bl[181] br[181] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_184 
+ bl[182] br[182] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_185 
+ bl[183] br[183] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_186 
+ bl[184] br[184] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_187 
+ bl[185] br[185] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_188 
+ bl[186] br[186] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_189 
+ bl[187] br[187] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_190 
+ bl[188] br[188] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_191 
+ bl[189] br[189] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_192 
+ bl[190] br[190] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_193 
+ bl[191] br[191] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_194 
+ bl[192] br[192] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_195 
+ bl[193] br[193] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_196 
+ bl[194] br[194] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_197 
+ bl[195] br[195] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_198 
+ bl[196] br[196] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_199 
+ bl[197] br[197] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_200 
+ bl[198] br[198] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_201 
+ bl[199] br[199] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_202 
+ bl[200] br[200] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_203 
+ bl[201] br[201] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_204 
+ bl[202] br[202] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_205 
+ bl[203] br[203] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_206 
+ bl[204] br[204] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_207 
+ bl[205] br[205] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_208 
+ bl[206] br[206] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_209 
+ bl[207] br[207] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_210 
+ bl[208] br[208] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_211 
+ bl[209] br[209] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_212 
+ bl[210] br[210] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_213 
+ bl[211] br[211] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_214 
+ bl[212] br[212] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_215 
+ bl[213] br[213] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_216 
+ bl[214] br[214] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_217 
+ bl[215] br[215] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_218 
+ bl[216] br[216] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_219 
+ bl[217] br[217] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_220 
+ bl[218] br[218] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_221 
+ bl[219] br[219] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_222 
+ bl[220] br[220] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_223 
+ bl[221] br[221] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_224 
+ bl[222] br[222] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_225 
+ bl[223] br[223] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_226 
+ bl[224] br[224] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_227 
+ bl[225] br[225] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_228 
+ bl[226] br[226] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_229 
+ bl[227] br[227] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_230 
+ bl[228] br[228] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_231 
+ bl[229] br[229] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_232 
+ bl[230] br[230] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_233 
+ bl[231] br[231] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_234 
+ bl[232] br[232] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_235 
+ bl[233] br[233] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_236 
+ bl[234] br[234] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_237 
+ bl[235] br[235] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_238 
+ bl[236] br[236] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_239 
+ bl[237] br[237] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_240 
+ bl[238] br[238] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_241 
+ bl[239] br[239] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_242 
+ bl[240] br[240] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_243 
+ bl[241] br[241] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_244 
+ bl[242] br[242] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_245 
+ bl[243] br[243] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_246 
+ bl[244] br[244] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_247 
+ bl[245] br[245] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_248 
+ bl[246] br[246] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_249 
+ bl[247] br[247] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_250 
+ bl[248] br[248] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_251 
+ bl[249] br[249] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_252 
+ bl[250] br[250] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_253 
+ bl[251] br[251] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_254 
+ bl[252] br[252] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_255 
+ bl[253] br[253] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_256 
+ bl[254] br[254] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_257 
+ bl[255] br[255] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_258 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_259 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_0 
+ vdd vdd vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_1 
+ rbl rbr vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_2 
+ bl[0] br[0] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_3 
+ bl[1] br[1] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_4 
+ bl[2] br[2] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_5 
+ bl[3] br[3] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_6 
+ bl[4] br[4] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_7 
+ bl[5] br[5] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_8 
+ bl[6] br[6] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_9 
+ bl[7] br[7] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_10 
+ bl[8] br[8] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_11 
+ bl[9] br[9] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_12 
+ bl[10] br[10] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_13 
+ bl[11] br[11] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_14 
+ bl[12] br[12] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_15 
+ bl[13] br[13] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_16 
+ bl[14] br[14] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_17 
+ bl[15] br[15] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_18 
+ bl[16] br[16] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_19 
+ bl[17] br[17] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_20 
+ bl[18] br[18] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_21 
+ bl[19] br[19] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_22 
+ bl[20] br[20] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_23 
+ bl[21] br[21] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_24 
+ bl[22] br[22] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_25 
+ bl[23] br[23] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_26 
+ bl[24] br[24] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_27 
+ bl[25] br[25] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_28 
+ bl[26] br[26] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_29 
+ bl[27] br[27] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_30 
+ bl[28] br[28] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_31 
+ bl[29] br[29] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_32 
+ bl[30] br[30] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_33 
+ bl[31] br[31] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_34 
+ bl[32] br[32] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_35 
+ bl[33] br[33] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_36 
+ bl[34] br[34] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_37 
+ bl[35] br[35] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_38 
+ bl[36] br[36] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_39 
+ bl[37] br[37] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_40 
+ bl[38] br[38] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_41 
+ bl[39] br[39] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_42 
+ bl[40] br[40] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_43 
+ bl[41] br[41] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_44 
+ bl[42] br[42] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_45 
+ bl[43] br[43] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_46 
+ bl[44] br[44] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_47 
+ bl[45] br[45] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_48 
+ bl[46] br[46] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_49 
+ bl[47] br[47] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_50 
+ bl[48] br[48] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_51 
+ bl[49] br[49] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_52 
+ bl[50] br[50] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_53 
+ bl[51] br[51] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_54 
+ bl[52] br[52] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_55 
+ bl[53] br[53] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_56 
+ bl[54] br[54] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_57 
+ bl[55] br[55] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_58 
+ bl[56] br[56] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_59 
+ bl[57] br[57] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_60 
+ bl[58] br[58] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_61 
+ bl[59] br[59] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_62 
+ bl[60] br[60] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_63 
+ bl[61] br[61] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_64 
+ bl[62] br[62] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_65 
+ bl[63] br[63] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_66 
+ bl[64] br[64] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_67 
+ bl[65] br[65] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_68 
+ bl[66] br[66] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_69 
+ bl[67] br[67] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_70 
+ bl[68] br[68] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_71 
+ bl[69] br[69] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_72 
+ bl[70] br[70] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_73 
+ bl[71] br[71] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_74 
+ bl[72] br[72] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_75 
+ bl[73] br[73] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_76 
+ bl[74] br[74] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_77 
+ bl[75] br[75] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_78 
+ bl[76] br[76] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_79 
+ bl[77] br[77] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_80 
+ bl[78] br[78] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_81 
+ bl[79] br[79] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_82 
+ bl[80] br[80] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_83 
+ bl[81] br[81] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_84 
+ bl[82] br[82] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_85 
+ bl[83] br[83] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_86 
+ bl[84] br[84] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_87 
+ bl[85] br[85] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_88 
+ bl[86] br[86] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_89 
+ bl[87] br[87] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_90 
+ bl[88] br[88] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_91 
+ bl[89] br[89] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_92 
+ bl[90] br[90] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_93 
+ bl[91] br[91] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_94 
+ bl[92] br[92] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_95 
+ bl[93] br[93] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_96 
+ bl[94] br[94] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_97 
+ bl[95] br[95] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_98 
+ bl[96] br[96] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_99 
+ bl[97] br[97] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_100 
+ bl[98] br[98] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_101 
+ bl[99] br[99] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_102 
+ bl[100] br[100] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_103 
+ bl[101] br[101] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_104 
+ bl[102] br[102] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_105 
+ bl[103] br[103] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_106 
+ bl[104] br[104] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_107 
+ bl[105] br[105] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_108 
+ bl[106] br[106] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_109 
+ bl[107] br[107] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_110 
+ bl[108] br[108] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_111 
+ bl[109] br[109] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_112 
+ bl[110] br[110] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_113 
+ bl[111] br[111] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_114 
+ bl[112] br[112] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_115 
+ bl[113] br[113] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_116 
+ bl[114] br[114] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_117 
+ bl[115] br[115] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_118 
+ bl[116] br[116] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_119 
+ bl[117] br[117] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_120 
+ bl[118] br[118] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_121 
+ bl[119] br[119] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_122 
+ bl[120] br[120] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_123 
+ bl[121] br[121] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_124 
+ bl[122] br[122] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_125 
+ bl[123] br[123] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_126 
+ bl[124] br[124] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_127 
+ bl[125] br[125] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_128 
+ bl[126] br[126] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_129 
+ bl[127] br[127] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_130 
+ bl[128] br[128] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_131 
+ bl[129] br[129] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_132 
+ bl[130] br[130] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_133 
+ bl[131] br[131] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_134 
+ bl[132] br[132] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_135 
+ bl[133] br[133] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_136 
+ bl[134] br[134] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_137 
+ bl[135] br[135] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_138 
+ bl[136] br[136] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_139 
+ bl[137] br[137] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_140 
+ bl[138] br[138] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_141 
+ bl[139] br[139] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_142 
+ bl[140] br[140] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_143 
+ bl[141] br[141] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_144 
+ bl[142] br[142] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_145 
+ bl[143] br[143] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_146 
+ bl[144] br[144] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_147 
+ bl[145] br[145] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_148 
+ bl[146] br[146] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_149 
+ bl[147] br[147] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_150 
+ bl[148] br[148] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_151 
+ bl[149] br[149] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_152 
+ bl[150] br[150] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_153 
+ bl[151] br[151] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_154 
+ bl[152] br[152] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_155 
+ bl[153] br[153] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_156 
+ bl[154] br[154] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_157 
+ bl[155] br[155] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_158 
+ bl[156] br[156] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_159 
+ bl[157] br[157] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_160 
+ bl[158] br[158] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_161 
+ bl[159] br[159] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_162 
+ bl[160] br[160] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_163 
+ bl[161] br[161] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_164 
+ bl[162] br[162] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_165 
+ bl[163] br[163] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_166 
+ bl[164] br[164] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_167 
+ bl[165] br[165] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_168 
+ bl[166] br[166] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_169 
+ bl[167] br[167] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_170 
+ bl[168] br[168] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_171 
+ bl[169] br[169] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_172 
+ bl[170] br[170] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_173 
+ bl[171] br[171] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_174 
+ bl[172] br[172] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_175 
+ bl[173] br[173] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_176 
+ bl[174] br[174] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_177 
+ bl[175] br[175] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_178 
+ bl[176] br[176] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_179 
+ bl[177] br[177] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_180 
+ bl[178] br[178] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_181 
+ bl[179] br[179] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_182 
+ bl[180] br[180] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_183 
+ bl[181] br[181] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_184 
+ bl[182] br[182] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_185 
+ bl[183] br[183] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_186 
+ bl[184] br[184] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_187 
+ bl[185] br[185] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_188 
+ bl[186] br[186] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_189 
+ bl[187] br[187] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_190 
+ bl[188] br[188] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_191 
+ bl[189] br[189] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_192 
+ bl[190] br[190] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_193 
+ bl[191] br[191] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_194 
+ bl[192] br[192] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_195 
+ bl[193] br[193] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_196 
+ bl[194] br[194] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_197 
+ bl[195] br[195] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_198 
+ bl[196] br[196] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_199 
+ bl[197] br[197] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_200 
+ bl[198] br[198] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_201 
+ bl[199] br[199] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_202 
+ bl[200] br[200] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_203 
+ bl[201] br[201] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_204 
+ bl[202] br[202] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_205 
+ bl[203] br[203] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_206 
+ bl[204] br[204] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_207 
+ bl[205] br[205] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_208 
+ bl[206] br[206] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_209 
+ bl[207] br[207] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_210 
+ bl[208] br[208] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_211 
+ bl[209] br[209] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_212 
+ bl[210] br[210] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_213 
+ bl[211] br[211] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_214 
+ bl[212] br[212] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_215 
+ bl[213] br[213] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_216 
+ bl[214] br[214] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_217 
+ bl[215] br[215] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_218 
+ bl[216] br[216] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_219 
+ bl[217] br[217] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_220 
+ bl[218] br[218] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_221 
+ bl[219] br[219] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_222 
+ bl[220] br[220] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_223 
+ bl[221] br[221] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_224 
+ bl[222] br[222] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_225 
+ bl[223] br[223] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_226 
+ bl[224] br[224] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_227 
+ bl[225] br[225] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_228 
+ bl[226] br[226] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_229 
+ bl[227] br[227] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_230 
+ bl[228] br[228] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_231 
+ bl[229] br[229] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_232 
+ bl[230] br[230] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_233 
+ bl[231] br[231] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_234 
+ bl[232] br[232] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_235 
+ bl[233] br[233] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_236 
+ bl[234] br[234] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_237 
+ bl[235] br[235] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_238 
+ bl[236] br[236] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_239 
+ bl[237] br[237] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_240 
+ bl[238] br[238] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_241 
+ bl[239] br[239] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_242 
+ bl[240] br[240] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_243 
+ bl[241] br[241] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_244 
+ bl[242] br[242] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_245 
+ bl[243] br[243] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_246 
+ bl[244] br[244] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_247 
+ bl[245] br[245] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_248 
+ bl[246] br[246] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_249 
+ bl[247] br[247] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_250 
+ bl[248] br[248] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_251 
+ bl[249] br[249] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_252 
+ bl[250] br[250] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_253 
+ bl[251] br[251] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_254 
+ bl[252] br[252] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_255 
+ bl[253] br[253] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_256 
+ bl[254] br[254] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_257 
+ bl[255] br[255] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_258 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_259 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_0 
+ vdd vdd vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_1 
+ rbl rbr vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_2 
+ bl[0] br[0] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_3 
+ bl[1] br[1] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_4 
+ bl[2] br[2] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_5 
+ bl[3] br[3] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_6 
+ bl[4] br[4] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_7 
+ bl[5] br[5] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_8 
+ bl[6] br[6] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_9 
+ bl[7] br[7] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_10 
+ bl[8] br[8] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_11 
+ bl[9] br[9] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_12 
+ bl[10] br[10] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_13 
+ bl[11] br[11] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_14 
+ bl[12] br[12] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_15 
+ bl[13] br[13] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_16 
+ bl[14] br[14] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_17 
+ bl[15] br[15] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_18 
+ bl[16] br[16] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_19 
+ bl[17] br[17] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_20 
+ bl[18] br[18] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_21 
+ bl[19] br[19] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_22 
+ bl[20] br[20] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_23 
+ bl[21] br[21] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_24 
+ bl[22] br[22] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_25 
+ bl[23] br[23] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_26 
+ bl[24] br[24] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_27 
+ bl[25] br[25] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_28 
+ bl[26] br[26] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_29 
+ bl[27] br[27] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_30 
+ bl[28] br[28] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_31 
+ bl[29] br[29] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_32 
+ bl[30] br[30] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_33 
+ bl[31] br[31] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_34 
+ bl[32] br[32] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_35 
+ bl[33] br[33] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_36 
+ bl[34] br[34] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_37 
+ bl[35] br[35] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_38 
+ bl[36] br[36] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_39 
+ bl[37] br[37] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_40 
+ bl[38] br[38] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_41 
+ bl[39] br[39] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_42 
+ bl[40] br[40] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_43 
+ bl[41] br[41] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_44 
+ bl[42] br[42] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_45 
+ bl[43] br[43] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_46 
+ bl[44] br[44] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_47 
+ bl[45] br[45] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_48 
+ bl[46] br[46] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_49 
+ bl[47] br[47] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_50 
+ bl[48] br[48] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_51 
+ bl[49] br[49] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_52 
+ bl[50] br[50] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_53 
+ bl[51] br[51] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_54 
+ bl[52] br[52] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_55 
+ bl[53] br[53] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_56 
+ bl[54] br[54] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_57 
+ bl[55] br[55] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_58 
+ bl[56] br[56] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_59 
+ bl[57] br[57] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_60 
+ bl[58] br[58] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_61 
+ bl[59] br[59] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_62 
+ bl[60] br[60] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_63 
+ bl[61] br[61] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_64 
+ bl[62] br[62] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_65 
+ bl[63] br[63] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_66 
+ bl[64] br[64] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_67 
+ bl[65] br[65] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_68 
+ bl[66] br[66] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_69 
+ bl[67] br[67] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_70 
+ bl[68] br[68] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_71 
+ bl[69] br[69] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_72 
+ bl[70] br[70] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_73 
+ bl[71] br[71] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_74 
+ bl[72] br[72] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_75 
+ bl[73] br[73] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_76 
+ bl[74] br[74] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_77 
+ bl[75] br[75] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_78 
+ bl[76] br[76] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_79 
+ bl[77] br[77] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_80 
+ bl[78] br[78] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_81 
+ bl[79] br[79] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_82 
+ bl[80] br[80] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_83 
+ bl[81] br[81] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_84 
+ bl[82] br[82] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_85 
+ bl[83] br[83] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_86 
+ bl[84] br[84] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_87 
+ bl[85] br[85] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_88 
+ bl[86] br[86] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_89 
+ bl[87] br[87] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_90 
+ bl[88] br[88] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_91 
+ bl[89] br[89] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_92 
+ bl[90] br[90] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_93 
+ bl[91] br[91] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_94 
+ bl[92] br[92] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_95 
+ bl[93] br[93] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_96 
+ bl[94] br[94] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_97 
+ bl[95] br[95] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_98 
+ bl[96] br[96] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_99 
+ bl[97] br[97] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_100 
+ bl[98] br[98] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_101 
+ bl[99] br[99] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_102 
+ bl[100] br[100] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_103 
+ bl[101] br[101] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_104 
+ bl[102] br[102] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_105 
+ bl[103] br[103] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_106 
+ bl[104] br[104] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_107 
+ bl[105] br[105] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_108 
+ bl[106] br[106] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_109 
+ bl[107] br[107] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_110 
+ bl[108] br[108] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_111 
+ bl[109] br[109] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_112 
+ bl[110] br[110] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_113 
+ bl[111] br[111] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_114 
+ bl[112] br[112] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_115 
+ bl[113] br[113] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_116 
+ bl[114] br[114] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_117 
+ bl[115] br[115] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_118 
+ bl[116] br[116] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_119 
+ bl[117] br[117] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_120 
+ bl[118] br[118] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_121 
+ bl[119] br[119] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_122 
+ bl[120] br[120] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_123 
+ bl[121] br[121] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_124 
+ bl[122] br[122] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_125 
+ bl[123] br[123] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_126 
+ bl[124] br[124] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_127 
+ bl[125] br[125] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_128 
+ bl[126] br[126] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_129 
+ bl[127] br[127] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_130 
+ bl[128] br[128] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_131 
+ bl[129] br[129] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_132 
+ bl[130] br[130] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_133 
+ bl[131] br[131] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_134 
+ bl[132] br[132] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_135 
+ bl[133] br[133] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_136 
+ bl[134] br[134] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_137 
+ bl[135] br[135] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_138 
+ bl[136] br[136] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_139 
+ bl[137] br[137] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_140 
+ bl[138] br[138] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_141 
+ bl[139] br[139] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_142 
+ bl[140] br[140] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_143 
+ bl[141] br[141] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_144 
+ bl[142] br[142] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_145 
+ bl[143] br[143] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_146 
+ bl[144] br[144] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_147 
+ bl[145] br[145] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_148 
+ bl[146] br[146] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_149 
+ bl[147] br[147] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_150 
+ bl[148] br[148] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_151 
+ bl[149] br[149] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_152 
+ bl[150] br[150] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_153 
+ bl[151] br[151] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_154 
+ bl[152] br[152] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_155 
+ bl[153] br[153] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_156 
+ bl[154] br[154] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_157 
+ bl[155] br[155] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_158 
+ bl[156] br[156] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_159 
+ bl[157] br[157] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_160 
+ bl[158] br[158] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_161 
+ bl[159] br[159] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_162 
+ bl[160] br[160] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_163 
+ bl[161] br[161] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_164 
+ bl[162] br[162] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_165 
+ bl[163] br[163] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_166 
+ bl[164] br[164] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_167 
+ bl[165] br[165] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_168 
+ bl[166] br[166] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_169 
+ bl[167] br[167] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_170 
+ bl[168] br[168] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_171 
+ bl[169] br[169] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_172 
+ bl[170] br[170] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_173 
+ bl[171] br[171] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_174 
+ bl[172] br[172] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_175 
+ bl[173] br[173] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_176 
+ bl[174] br[174] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_177 
+ bl[175] br[175] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_178 
+ bl[176] br[176] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_179 
+ bl[177] br[177] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_180 
+ bl[178] br[178] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_181 
+ bl[179] br[179] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_182 
+ bl[180] br[180] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_183 
+ bl[181] br[181] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_184 
+ bl[182] br[182] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_185 
+ bl[183] br[183] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_186 
+ bl[184] br[184] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_187 
+ bl[185] br[185] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_188 
+ bl[186] br[186] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_189 
+ bl[187] br[187] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_190 
+ bl[188] br[188] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_191 
+ bl[189] br[189] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_192 
+ bl[190] br[190] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_193 
+ bl[191] br[191] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_194 
+ bl[192] br[192] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_195 
+ bl[193] br[193] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_196 
+ bl[194] br[194] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_197 
+ bl[195] br[195] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_198 
+ bl[196] br[196] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_199 
+ bl[197] br[197] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_200 
+ bl[198] br[198] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_201 
+ bl[199] br[199] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_202 
+ bl[200] br[200] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_203 
+ bl[201] br[201] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_204 
+ bl[202] br[202] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_205 
+ bl[203] br[203] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_206 
+ bl[204] br[204] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_207 
+ bl[205] br[205] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_208 
+ bl[206] br[206] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_209 
+ bl[207] br[207] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_210 
+ bl[208] br[208] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_211 
+ bl[209] br[209] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_212 
+ bl[210] br[210] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_213 
+ bl[211] br[211] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_214 
+ bl[212] br[212] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_215 
+ bl[213] br[213] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_216 
+ bl[214] br[214] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_217 
+ bl[215] br[215] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_218 
+ bl[216] br[216] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_219 
+ bl[217] br[217] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_220 
+ bl[218] br[218] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_221 
+ bl[219] br[219] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_222 
+ bl[220] br[220] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_223 
+ bl[221] br[221] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_224 
+ bl[222] br[222] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_225 
+ bl[223] br[223] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_226 
+ bl[224] br[224] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_227 
+ bl[225] br[225] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_228 
+ bl[226] br[226] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_229 
+ bl[227] br[227] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_230 
+ bl[228] br[228] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_231 
+ bl[229] br[229] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_232 
+ bl[230] br[230] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_233 
+ bl[231] br[231] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_234 
+ bl[232] br[232] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_235 
+ bl[233] br[233] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_236 
+ bl[234] br[234] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_237 
+ bl[235] br[235] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_238 
+ bl[236] br[236] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_239 
+ bl[237] br[237] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_240 
+ bl[238] br[238] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_241 
+ bl[239] br[239] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_242 
+ bl[240] br[240] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_243 
+ bl[241] br[241] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_244 
+ bl[242] br[242] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_245 
+ bl[243] br[243] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_246 
+ bl[244] br[244] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_247 
+ bl[245] br[245] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_248 
+ bl[246] br[246] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_249 
+ bl[247] br[247] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_250 
+ bl[248] br[248] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_251 
+ bl[249] br[249] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_252 
+ bl[250] br[250] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_253 
+ bl[251] br[251] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_254 
+ bl[252] br[252] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_255 
+ bl[253] br[253] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_256 
+ bl[254] br[254] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_257 
+ bl[255] br[255] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_258 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_259 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xcolend_0_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_0_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_bot 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_top 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_bot 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_top 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_bot 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_top 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_bot 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_top 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_bot 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_top 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_bot 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_top 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_bot 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_top 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_bot 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_top 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_bot 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_top 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_bot 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_top 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_bot 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_top 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_bot 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_top 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_bot 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_top 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_bot 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_top 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_bot 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_top 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_bot 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_top 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_bot 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_top 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_bot 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_top 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_bot 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_top 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_bot 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_top 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_bot 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_top 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_bot 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_top 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_bot 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_top 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_bot 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_top 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_bot 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_top 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_bot 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_top 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_bot 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_top 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_bot 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_top 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_bot 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_top 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_bot 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_top 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_bot 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_top 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_bot 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_top 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_bot 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_top 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_bot 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_top 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_bot 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_top 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_bot 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_top 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_bot 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_top 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_bot 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_top 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_bot 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_top 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_bot 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_top 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_bot 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_top 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_bot 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_top 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_bot 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_top 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_bot 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_top 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_bot 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_top 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_bot 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_top 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_bot 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_top 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_bot 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_top 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_bot 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_top 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_bot 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_top 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_bot 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_top 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_bot 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_top 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_bot 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_top 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_bot 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_top 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_bot 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_top 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_bot 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_top 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_bot 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_top 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_bot 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_top 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_bot 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_top 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_bot 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_top 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_bot 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_top 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_bot 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_top 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_bot 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_top 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_bot 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_top 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_bot 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_top 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_bot 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_top 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_bot 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_top 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_bot 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_top 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_bot 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_top 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_bot 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_top 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_bot 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_top 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_bot 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_top 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_bot 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_top 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_bot 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_top 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_bot 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_top 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_bot 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_top 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_bot 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_top 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_bot 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_top 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_bot 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_top 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_bot 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_top 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_bot 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_top 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_bot 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_top 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_bot 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_top 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_bot 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_top 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_bot 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_top 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_bot 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_top 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_bot 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_top 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_bot 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_top 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_bot 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_top 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_bot 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_top 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_bot 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_top 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_bot 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_top 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_bot 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_top 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_bot 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_top 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_bot 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_top 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_bot 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_top 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_bot 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_top 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_bot 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_top 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_bot 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_top 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_bot 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_top 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_bot 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_top 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_bot 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_top 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_bot 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_top 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_bot 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_top 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_bot 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_top 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_bot 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_top 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_bot 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_top 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_bot 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_top 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_bot 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_top 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_bot 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_top 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_bot 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_top 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_bot 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_top 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_bot 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_top 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_bot 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_top 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_bot 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_top 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_bot 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_top 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_bot 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_top 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_bot 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_top 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_bot 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_top 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_bot 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_top 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_bot 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_top 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_bot 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_top 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_bot 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_top 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_bot 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_top 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_bot 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_top 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_bot 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_top 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_bot 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_top 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_bot 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_top 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_bot 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_top 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_bot 
+ br[128] vdd vss bl[128] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_top 
+ br[128] vdd vss bl[128] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_bot 
+ br[129] vdd vss bl[129] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_top 
+ br[129] vdd vss bl[129] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_132_bot 
+ br[130] vdd vss bl[130] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_132_top 
+ br[130] vdd vss bl[130] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_133_bot 
+ br[131] vdd vss bl[131] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_133_top 
+ br[131] vdd vss bl[131] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_134_bot 
+ br[132] vdd vss bl[132] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_134_top 
+ br[132] vdd vss bl[132] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_135_bot 
+ br[133] vdd vss bl[133] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_135_top 
+ br[133] vdd vss bl[133] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_136_bot 
+ br[134] vdd vss bl[134] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_136_top 
+ br[134] vdd vss bl[134] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_137_bot 
+ br[135] vdd vss bl[135] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_137_top 
+ br[135] vdd vss bl[135] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_138_bot 
+ br[136] vdd vss bl[136] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_138_top 
+ br[136] vdd vss bl[136] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_139_bot 
+ br[137] vdd vss bl[137] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_139_top 
+ br[137] vdd vss bl[137] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_140_bot 
+ br[138] vdd vss bl[138] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_140_top 
+ br[138] vdd vss bl[138] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_141_bot 
+ br[139] vdd vss bl[139] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_141_top 
+ br[139] vdd vss bl[139] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_142_bot 
+ br[140] vdd vss bl[140] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_142_top 
+ br[140] vdd vss bl[140] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_143_bot 
+ br[141] vdd vss bl[141] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_143_top 
+ br[141] vdd vss bl[141] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_144_bot 
+ br[142] vdd vss bl[142] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_144_top 
+ br[142] vdd vss bl[142] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_145_bot 
+ br[143] vdd vss bl[143] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_145_top 
+ br[143] vdd vss bl[143] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_146_bot 
+ br[144] vdd vss bl[144] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_146_top 
+ br[144] vdd vss bl[144] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_147_bot 
+ br[145] vdd vss bl[145] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_147_top 
+ br[145] vdd vss bl[145] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_148_bot 
+ br[146] vdd vss bl[146] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_148_top 
+ br[146] vdd vss bl[146] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_149_bot 
+ br[147] vdd vss bl[147] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_149_top 
+ br[147] vdd vss bl[147] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_150_bot 
+ br[148] vdd vss bl[148] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_150_top 
+ br[148] vdd vss bl[148] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_151_bot 
+ br[149] vdd vss bl[149] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_151_top 
+ br[149] vdd vss bl[149] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_152_bot 
+ br[150] vdd vss bl[150] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_152_top 
+ br[150] vdd vss bl[150] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_153_bot 
+ br[151] vdd vss bl[151] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_153_top 
+ br[151] vdd vss bl[151] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_154_bot 
+ br[152] vdd vss bl[152] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_154_top 
+ br[152] vdd vss bl[152] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_155_bot 
+ br[153] vdd vss bl[153] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_155_top 
+ br[153] vdd vss bl[153] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_156_bot 
+ br[154] vdd vss bl[154] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_156_top 
+ br[154] vdd vss bl[154] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_157_bot 
+ br[155] vdd vss bl[155] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_157_top 
+ br[155] vdd vss bl[155] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_158_bot 
+ br[156] vdd vss bl[156] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_158_top 
+ br[156] vdd vss bl[156] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_159_bot 
+ br[157] vdd vss bl[157] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_159_top 
+ br[157] vdd vss bl[157] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_160_bot 
+ br[158] vdd vss bl[158] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_160_top 
+ br[158] vdd vss bl[158] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_161_bot 
+ br[159] vdd vss bl[159] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_161_top 
+ br[159] vdd vss bl[159] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_162_bot 
+ br[160] vdd vss bl[160] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_162_top 
+ br[160] vdd vss bl[160] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_163_bot 
+ br[161] vdd vss bl[161] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_163_top 
+ br[161] vdd vss bl[161] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_164_bot 
+ br[162] vdd vss bl[162] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_164_top 
+ br[162] vdd vss bl[162] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_165_bot 
+ br[163] vdd vss bl[163] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_165_top 
+ br[163] vdd vss bl[163] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_166_bot 
+ br[164] vdd vss bl[164] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_166_top 
+ br[164] vdd vss bl[164] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_167_bot 
+ br[165] vdd vss bl[165] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_167_top 
+ br[165] vdd vss bl[165] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_168_bot 
+ br[166] vdd vss bl[166] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_168_top 
+ br[166] vdd vss bl[166] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_169_bot 
+ br[167] vdd vss bl[167] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_169_top 
+ br[167] vdd vss bl[167] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_170_bot 
+ br[168] vdd vss bl[168] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_170_top 
+ br[168] vdd vss bl[168] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_171_bot 
+ br[169] vdd vss bl[169] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_171_top 
+ br[169] vdd vss bl[169] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_172_bot 
+ br[170] vdd vss bl[170] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_172_top 
+ br[170] vdd vss bl[170] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_173_bot 
+ br[171] vdd vss bl[171] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_173_top 
+ br[171] vdd vss bl[171] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_174_bot 
+ br[172] vdd vss bl[172] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_174_top 
+ br[172] vdd vss bl[172] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_175_bot 
+ br[173] vdd vss bl[173] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_175_top 
+ br[173] vdd vss bl[173] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_176_bot 
+ br[174] vdd vss bl[174] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_176_top 
+ br[174] vdd vss bl[174] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_177_bot 
+ br[175] vdd vss bl[175] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_177_top 
+ br[175] vdd vss bl[175] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_178_bot 
+ br[176] vdd vss bl[176] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_178_top 
+ br[176] vdd vss bl[176] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_179_bot 
+ br[177] vdd vss bl[177] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_179_top 
+ br[177] vdd vss bl[177] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_180_bot 
+ br[178] vdd vss bl[178] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_180_top 
+ br[178] vdd vss bl[178] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_181_bot 
+ br[179] vdd vss bl[179] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_181_top 
+ br[179] vdd vss bl[179] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_182_bot 
+ br[180] vdd vss bl[180] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_182_top 
+ br[180] vdd vss bl[180] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_183_bot 
+ br[181] vdd vss bl[181] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_183_top 
+ br[181] vdd vss bl[181] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_184_bot 
+ br[182] vdd vss bl[182] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_184_top 
+ br[182] vdd vss bl[182] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_185_bot 
+ br[183] vdd vss bl[183] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_185_top 
+ br[183] vdd vss bl[183] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_186_bot 
+ br[184] vdd vss bl[184] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_186_top 
+ br[184] vdd vss bl[184] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_187_bot 
+ br[185] vdd vss bl[185] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_187_top 
+ br[185] vdd vss bl[185] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_188_bot 
+ br[186] vdd vss bl[186] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_188_top 
+ br[186] vdd vss bl[186] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_189_bot 
+ br[187] vdd vss bl[187] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_189_top 
+ br[187] vdd vss bl[187] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_190_bot 
+ br[188] vdd vss bl[188] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_190_top 
+ br[188] vdd vss bl[188] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_191_bot 
+ br[189] vdd vss bl[189] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_191_top 
+ br[189] vdd vss bl[189] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_192_bot 
+ br[190] vdd vss bl[190] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_192_top 
+ br[190] vdd vss bl[190] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_193_bot 
+ br[191] vdd vss bl[191] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_193_top 
+ br[191] vdd vss bl[191] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_194_bot 
+ br[192] vdd vss bl[192] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_194_top 
+ br[192] vdd vss bl[192] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_195_bot 
+ br[193] vdd vss bl[193] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_195_top 
+ br[193] vdd vss bl[193] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_196_bot 
+ br[194] vdd vss bl[194] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_196_top 
+ br[194] vdd vss bl[194] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_197_bot 
+ br[195] vdd vss bl[195] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_197_top 
+ br[195] vdd vss bl[195] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_198_bot 
+ br[196] vdd vss bl[196] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_198_top 
+ br[196] vdd vss bl[196] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_199_bot 
+ br[197] vdd vss bl[197] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_199_top 
+ br[197] vdd vss bl[197] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_200_bot 
+ br[198] vdd vss bl[198] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_200_top 
+ br[198] vdd vss bl[198] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_201_bot 
+ br[199] vdd vss bl[199] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_201_top 
+ br[199] vdd vss bl[199] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_202_bot 
+ br[200] vdd vss bl[200] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_202_top 
+ br[200] vdd vss bl[200] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_203_bot 
+ br[201] vdd vss bl[201] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_203_top 
+ br[201] vdd vss bl[201] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_204_bot 
+ br[202] vdd vss bl[202] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_204_top 
+ br[202] vdd vss bl[202] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_205_bot 
+ br[203] vdd vss bl[203] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_205_top 
+ br[203] vdd vss bl[203] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_206_bot 
+ br[204] vdd vss bl[204] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_206_top 
+ br[204] vdd vss bl[204] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_207_bot 
+ br[205] vdd vss bl[205] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_207_top 
+ br[205] vdd vss bl[205] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_208_bot 
+ br[206] vdd vss bl[206] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_208_top 
+ br[206] vdd vss bl[206] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_209_bot 
+ br[207] vdd vss bl[207] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_209_top 
+ br[207] vdd vss bl[207] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_210_bot 
+ br[208] vdd vss bl[208] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_210_top 
+ br[208] vdd vss bl[208] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_211_bot 
+ br[209] vdd vss bl[209] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_211_top 
+ br[209] vdd vss bl[209] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_212_bot 
+ br[210] vdd vss bl[210] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_212_top 
+ br[210] vdd vss bl[210] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_213_bot 
+ br[211] vdd vss bl[211] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_213_top 
+ br[211] vdd vss bl[211] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_214_bot 
+ br[212] vdd vss bl[212] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_214_top 
+ br[212] vdd vss bl[212] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_215_bot 
+ br[213] vdd vss bl[213] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_215_top 
+ br[213] vdd vss bl[213] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_216_bot 
+ br[214] vdd vss bl[214] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_216_top 
+ br[214] vdd vss bl[214] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_217_bot 
+ br[215] vdd vss bl[215] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_217_top 
+ br[215] vdd vss bl[215] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_218_bot 
+ br[216] vdd vss bl[216] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_218_top 
+ br[216] vdd vss bl[216] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_219_bot 
+ br[217] vdd vss bl[217] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_219_top 
+ br[217] vdd vss bl[217] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_220_bot 
+ br[218] vdd vss bl[218] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_220_top 
+ br[218] vdd vss bl[218] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_221_bot 
+ br[219] vdd vss bl[219] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_221_top 
+ br[219] vdd vss bl[219] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_222_bot 
+ br[220] vdd vss bl[220] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_222_top 
+ br[220] vdd vss bl[220] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_223_bot 
+ br[221] vdd vss bl[221] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_223_top 
+ br[221] vdd vss bl[221] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_224_bot 
+ br[222] vdd vss bl[222] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_224_top 
+ br[222] vdd vss bl[222] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_225_bot 
+ br[223] vdd vss bl[223] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_225_top 
+ br[223] vdd vss bl[223] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_226_bot 
+ br[224] vdd vss bl[224] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_226_top 
+ br[224] vdd vss bl[224] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_227_bot 
+ br[225] vdd vss bl[225] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_227_top 
+ br[225] vdd vss bl[225] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_228_bot 
+ br[226] vdd vss bl[226] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_228_top 
+ br[226] vdd vss bl[226] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_229_bot 
+ br[227] vdd vss bl[227] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_229_top 
+ br[227] vdd vss bl[227] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_230_bot 
+ br[228] vdd vss bl[228] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_230_top 
+ br[228] vdd vss bl[228] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_231_bot 
+ br[229] vdd vss bl[229] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_231_top 
+ br[229] vdd vss bl[229] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_232_bot 
+ br[230] vdd vss bl[230] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_232_top 
+ br[230] vdd vss bl[230] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_233_bot 
+ br[231] vdd vss bl[231] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_233_top 
+ br[231] vdd vss bl[231] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_234_bot 
+ br[232] vdd vss bl[232] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_234_top 
+ br[232] vdd vss bl[232] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_235_bot 
+ br[233] vdd vss bl[233] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_235_top 
+ br[233] vdd vss bl[233] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_236_bot 
+ br[234] vdd vss bl[234] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_236_top 
+ br[234] vdd vss bl[234] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_237_bot 
+ br[235] vdd vss bl[235] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_237_top 
+ br[235] vdd vss bl[235] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_238_bot 
+ br[236] vdd vss bl[236] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_238_top 
+ br[236] vdd vss bl[236] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_239_bot 
+ br[237] vdd vss bl[237] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_239_top 
+ br[237] vdd vss bl[237] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_240_bot 
+ br[238] vdd vss bl[238] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_240_top 
+ br[238] vdd vss bl[238] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_241_bot 
+ br[239] vdd vss bl[239] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_241_top 
+ br[239] vdd vss bl[239] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_242_bot 
+ br[240] vdd vss bl[240] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_242_top 
+ br[240] vdd vss bl[240] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_243_bot 
+ br[241] vdd vss bl[241] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_243_top 
+ br[241] vdd vss bl[241] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_244_bot 
+ br[242] vdd vss bl[242] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_244_top 
+ br[242] vdd vss bl[242] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_245_bot 
+ br[243] vdd vss bl[243] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_245_top 
+ br[243] vdd vss bl[243] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_246_bot 
+ br[244] vdd vss bl[244] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_246_top 
+ br[244] vdd vss bl[244] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_247_bot 
+ br[245] vdd vss bl[245] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_247_top 
+ br[245] vdd vss bl[245] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_248_bot 
+ br[246] vdd vss bl[246] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_248_top 
+ br[246] vdd vss bl[246] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_249_bot 
+ br[247] vdd vss bl[247] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_249_top 
+ br[247] vdd vss bl[247] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_250_bot 
+ br[248] vdd vss bl[248] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_250_top 
+ br[248] vdd vss bl[248] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_251_bot 
+ br[249] vdd vss bl[249] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_251_top 
+ br[249] vdd vss bl[249] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_252_bot 
+ br[250] vdd vss bl[250] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_252_top 
+ br[250] vdd vss bl[250] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_253_bot 
+ br[251] vdd vss bl[251] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_253_top 
+ br[251] vdd vss bl[251] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_254_bot 
+ br[252] vdd vss bl[252] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_254_top 
+ br[252] vdd vss bl[252] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_255_bot 
+ br[253] vdd vss bl[253] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_255_top 
+ br[253] vdd vss bl[253] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_256_bot 
+ br[254] vdd vss bl[254] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_256_top 
+ br[254] vdd vss bl[254] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_257_bot 
+ br[255] vdd vss bl[255] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_257_top 
+ br[255] vdd vss bl[255] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_258_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_258_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_259_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_259_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

.ENDS

.SUBCKT precharge 
+ vdd bl br en_b 

xbl_pull_up 
+ bl en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xbr_pull_up 
+ br en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xequalizer 
+ bl en_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

.ENDS

.SUBCKT precharge_array 
+ vdd en_b bl[256] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[256] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] 

xprecharge_0 
+ vdd bl[0] br[0] en_b 
+ precharge 
* No parameters

xprecharge_1 
+ vdd bl[1] br[1] en_b 
+ precharge 
* No parameters

xprecharge_2 
+ vdd bl[2] br[2] en_b 
+ precharge 
* No parameters

xprecharge_3 
+ vdd bl[3] br[3] en_b 
+ precharge 
* No parameters

xprecharge_4 
+ vdd bl[4] br[4] en_b 
+ precharge 
* No parameters

xprecharge_5 
+ vdd bl[5] br[5] en_b 
+ precharge 
* No parameters

xprecharge_6 
+ vdd bl[6] br[6] en_b 
+ precharge 
* No parameters

xprecharge_7 
+ vdd bl[7] br[7] en_b 
+ precharge 
* No parameters

xprecharge_8 
+ vdd bl[8] br[8] en_b 
+ precharge 
* No parameters

xprecharge_9 
+ vdd bl[9] br[9] en_b 
+ precharge 
* No parameters

xprecharge_10 
+ vdd bl[10] br[10] en_b 
+ precharge 
* No parameters

xprecharge_11 
+ vdd bl[11] br[11] en_b 
+ precharge 
* No parameters

xprecharge_12 
+ vdd bl[12] br[12] en_b 
+ precharge 
* No parameters

xprecharge_13 
+ vdd bl[13] br[13] en_b 
+ precharge 
* No parameters

xprecharge_14 
+ vdd bl[14] br[14] en_b 
+ precharge 
* No parameters

xprecharge_15 
+ vdd bl[15] br[15] en_b 
+ precharge 
* No parameters

xprecharge_16 
+ vdd bl[16] br[16] en_b 
+ precharge 
* No parameters

xprecharge_17 
+ vdd bl[17] br[17] en_b 
+ precharge 
* No parameters

xprecharge_18 
+ vdd bl[18] br[18] en_b 
+ precharge 
* No parameters

xprecharge_19 
+ vdd bl[19] br[19] en_b 
+ precharge 
* No parameters

xprecharge_20 
+ vdd bl[20] br[20] en_b 
+ precharge 
* No parameters

xprecharge_21 
+ vdd bl[21] br[21] en_b 
+ precharge 
* No parameters

xprecharge_22 
+ vdd bl[22] br[22] en_b 
+ precharge 
* No parameters

xprecharge_23 
+ vdd bl[23] br[23] en_b 
+ precharge 
* No parameters

xprecharge_24 
+ vdd bl[24] br[24] en_b 
+ precharge 
* No parameters

xprecharge_25 
+ vdd bl[25] br[25] en_b 
+ precharge 
* No parameters

xprecharge_26 
+ vdd bl[26] br[26] en_b 
+ precharge 
* No parameters

xprecharge_27 
+ vdd bl[27] br[27] en_b 
+ precharge 
* No parameters

xprecharge_28 
+ vdd bl[28] br[28] en_b 
+ precharge 
* No parameters

xprecharge_29 
+ vdd bl[29] br[29] en_b 
+ precharge 
* No parameters

xprecharge_30 
+ vdd bl[30] br[30] en_b 
+ precharge 
* No parameters

xprecharge_31 
+ vdd bl[31] br[31] en_b 
+ precharge 
* No parameters

xprecharge_32 
+ vdd bl[32] br[32] en_b 
+ precharge 
* No parameters

xprecharge_33 
+ vdd bl[33] br[33] en_b 
+ precharge 
* No parameters

xprecharge_34 
+ vdd bl[34] br[34] en_b 
+ precharge 
* No parameters

xprecharge_35 
+ vdd bl[35] br[35] en_b 
+ precharge 
* No parameters

xprecharge_36 
+ vdd bl[36] br[36] en_b 
+ precharge 
* No parameters

xprecharge_37 
+ vdd bl[37] br[37] en_b 
+ precharge 
* No parameters

xprecharge_38 
+ vdd bl[38] br[38] en_b 
+ precharge 
* No parameters

xprecharge_39 
+ vdd bl[39] br[39] en_b 
+ precharge 
* No parameters

xprecharge_40 
+ vdd bl[40] br[40] en_b 
+ precharge 
* No parameters

xprecharge_41 
+ vdd bl[41] br[41] en_b 
+ precharge 
* No parameters

xprecharge_42 
+ vdd bl[42] br[42] en_b 
+ precharge 
* No parameters

xprecharge_43 
+ vdd bl[43] br[43] en_b 
+ precharge 
* No parameters

xprecharge_44 
+ vdd bl[44] br[44] en_b 
+ precharge 
* No parameters

xprecharge_45 
+ vdd bl[45] br[45] en_b 
+ precharge 
* No parameters

xprecharge_46 
+ vdd bl[46] br[46] en_b 
+ precharge 
* No parameters

xprecharge_47 
+ vdd bl[47] br[47] en_b 
+ precharge 
* No parameters

xprecharge_48 
+ vdd bl[48] br[48] en_b 
+ precharge 
* No parameters

xprecharge_49 
+ vdd bl[49] br[49] en_b 
+ precharge 
* No parameters

xprecharge_50 
+ vdd bl[50] br[50] en_b 
+ precharge 
* No parameters

xprecharge_51 
+ vdd bl[51] br[51] en_b 
+ precharge 
* No parameters

xprecharge_52 
+ vdd bl[52] br[52] en_b 
+ precharge 
* No parameters

xprecharge_53 
+ vdd bl[53] br[53] en_b 
+ precharge 
* No parameters

xprecharge_54 
+ vdd bl[54] br[54] en_b 
+ precharge 
* No parameters

xprecharge_55 
+ vdd bl[55] br[55] en_b 
+ precharge 
* No parameters

xprecharge_56 
+ vdd bl[56] br[56] en_b 
+ precharge 
* No parameters

xprecharge_57 
+ vdd bl[57] br[57] en_b 
+ precharge 
* No parameters

xprecharge_58 
+ vdd bl[58] br[58] en_b 
+ precharge 
* No parameters

xprecharge_59 
+ vdd bl[59] br[59] en_b 
+ precharge 
* No parameters

xprecharge_60 
+ vdd bl[60] br[60] en_b 
+ precharge 
* No parameters

xprecharge_61 
+ vdd bl[61] br[61] en_b 
+ precharge 
* No parameters

xprecharge_62 
+ vdd bl[62] br[62] en_b 
+ precharge 
* No parameters

xprecharge_63 
+ vdd bl[63] br[63] en_b 
+ precharge 
* No parameters

xprecharge_64 
+ vdd bl[64] br[64] en_b 
+ precharge 
* No parameters

xprecharge_65 
+ vdd bl[65] br[65] en_b 
+ precharge 
* No parameters

xprecharge_66 
+ vdd bl[66] br[66] en_b 
+ precharge 
* No parameters

xprecharge_67 
+ vdd bl[67] br[67] en_b 
+ precharge 
* No parameters

xprecharge_68 
+ vdd bl[68] br[68] en_b 
+ precharge 
* No parameters

xprecharge_69 
+ vdd bl[69] br[69] en_b 
+ precharge 
* No parameters

xprecharge_70 
+ vdd bl[70] br[70] en_b 
+ precharge 
* No parameters

xprecharge_71 
+ vdd bl[71] br[71] en_b 
+ precharge 
* No parameters

xprecharge_72 
+ vdd bl[72] br[72] en_b 
+ precharge 
* No parameters

xprecharge_73 
+ vdd bl[73] br[73] en_b 
+ precharge 
* No parameters

xprecharge_74 
+ vdd bl[74] br[74] en_b 
+ precharge 
* No parameters

xprecharge_75 
+ vdd bl[75] br[75] en_b 
+ precharge 
* No parameters

xprecharge_76 
+ vdd bl[76] br[76] en_b 
+ precharge 
* No parameters

xprecharge_77 
+ vdd bl[77] br[77] en_b 
+ precharge 
* No parameters

xprecharge_78 
+ vdd bl[78] br[78] en_b 
+ precharge 
* No parameters

xprecharge_79 
+ vdd bl[79] br[79] en_b 
+ precharge 
* No parameters

xprecharge_80 
+ vdd bl[80] br[80] en_b 
+ precharge 
* No parameters

xprecharge_81 
+ vdd bl[81] br[81] en_b 
+ precharge 
* No parameters

xprecharge_82 
+ vdd bl[82] br[82] en_b 
+ precharge 
* No parameters

xprecharge_83 
+ vdd bl[83] br[83] en_b 
+ precharge 
* No parameters

xprecharge_84 
+ vdd bl[84] br[84] en_b 
+ precharge 
* No parameters

xprecharge_85 
+ vdd bl[85] br[85] en_b 
+ precharge 
* No parameters

xprecharge_86 
+ vdd bl[86] br[86] en_b 
+ precharge 
* No parameters

xprecharge_87 
+ vdd bl[87] br[87] en_b 
+ precharge 
* No parameters

xprecharge_88 
+ vdd bl[88] br[88] en_b 
+ precharge 
* No parameters

xprecharge_89 
+ vdd bl[89] br[89] en_b 
+ precharge 
* No parameters

xprecharge_90 
+ vdd bl[90] br[90] en_b 
+ precharge 
* No parameters

xprecharge_91 
+ vdd bl[91] br[91] en_b 
+ precharge 
* No parameters

xprecharge_92 
+ vdd bl[92] br[92] en_b 
+ precharge 
* No parameters

xprecharge_93 
+ vdd bl[93] br[93] en_b 
+ precharge 
* No parameters

xprecharge_94 
+ vdd bl[94] br[94] en_b 
+ precharge 
* No parameters

xprecharge_95 
+ vdd bl[95] br[95] en_b 
+ precharge 
* No parameters

xprecharge_96 
+ vdd bl[96] br[96] en_b 
+ precharge 
* No parameters

xprecharge_97 
+ vdd bl[97] br[97] en_b 
+ precharge 
* No parameters

xprecharge_98 
+ vdd bl[98] br[98] en_b 
+ precharge 
* No parameters

xprecharge_99 
+ vdd bl[99] br[99] en_b 
+ precharge 
* No parameters

xprecharge_100 
+ vdd bl[100] br[100] en_b 
+ precharge 
* No parameters

xprecharge_101 
+ vdd bl[101] br[101] en_b 
+ precharge 
* No parameters

xprecharge_102 
+ vdd bl[102] br[102] en_b 
+ precharge 
* No parameters

xprecharge_103 
+ vdd bl[103] br[103] en_b 
+ precharge 
* No parameters

xprecharge_104 
+ vdd bl[104] br[104] en_b 
+ precharge 
* No parameters

xprecharge_105 
+ vdd bl[105] br[105] en_b 
+ precharge 
* No parameters

xprecharge_106 
+ vdd bl[106] br[106] en_b 
+ precharge 
* No parameters

xprecharge_107 
+ vdd bl[107] br[107] en_b 
+ precharge 
* No parameters

xprecharge_108 
+ vdd bl[108] br[108] en_b 
+ precharge 
* No parameters

xprecharge_109 
+ vdd bl[109] br[109] en_b 
+ precharge 
* No parameters

xprecharge_110 
+ vdd bl[110] br[110] en_b 
+ precharge 
* No parameters

xprecharge_111 
+ vdd bl[111] br[111] en_b 
+ precharge 
* No parameters

xprecharge_112 
+ vdd bl[112] br[112] en_b 
+ precharge 
* No parameters

xprecharge_113 
+ vdd bl[113] br[113] en_b 
+ precharge 
* No parameters

xprecharge_114 
+ vdd bl[114] br[114] en_b 
+ precharge 
* No parameters

xprecharge_115 
+ vdd bl[115] br[115] en_b 
+ precharge 
* No parameters

xprecharge_116 
+ vdd bl[116] br[116] en_b 
+ precharge 
* No parameters

xprecharge_117 
+ vdd bl[117] br[117] en_b 
+ precharge 
* No parameters

xprecharge_118 
+ vdd bl[118] br[118] en_b 
+ precharge 
* No parameters

xprecharge_119 
+ vdd bl[119] br[119] en_b 
+ precharge 
* No parameters

xprecharge_120 
+ vdd bl[120] br[120] en_b 
+ precharge 
* No parameters

xprecharge_121 
+ vdd bl[121] br[121] en_b 
+ precharge 
* No parameters

xprecharge_122 
+ vdd bl[122] br[122] en_b 
+ precharge 
* No parameters

xprecharge_123 
+ vdd bl[123] br[123] en_b 
+ precharge 
* No parameters

xprecharge_124 
+ vdd bl[124] br[124] en_b 
+ precharge 
* No parameters

xprecharge_125 
+ vdd bl[125] br[125] en_b 
+ precharge 
* No parameters

xprecharge_126 
+ vdd bl[126] br[126] en_b 
+ precharge 
* No parameters

xprecharge_127 
+ vdd bl[127] br[127] en_b 
+ precharge 
* No parameters

xprecharge_128 
+ vdd bl[128] br[128] en_b 
+ precharge 
* No parameters

xprecharge_129 
+ vdd bl[129] br[129] en_b 
+ precharge 
* No parameters

xprecharge_130 
+ vdd bl[130] br[130] en_b 
+ precharge 
* No parameters

xprecharge_131 
+ vdd bl[131] br[131] en_b 
+ precharge 
* No parameters

xprecharge_132 
+ vdd bl[132] br[132] en_b 
+ precharge 
* No parameters

xprecharge_133 
+ vdd bl[133] br[133] en_b 
+ precharge 
* No parameters

xprecharge_134 
+ vdd bl[134] br[134] en_b 
+ precharge 
* No parameters

xprecharge_135 
+ vdd bl[135] br[135] en_b 
+ precharge 
* No parameters

xprecharge_136 
+ vdd bl[136] br[136] en_b 
+ precharge 
* No parameters

xprecharge_137 
+ vdd bl[137] br[137] en_b 
+ precharge 
* No parameters

xprecharge_138 
+ vdd bl[138] br[138] en_b 
+ precharge 
* No parameters

xprecharge_139 
+ vdd bl[139] br[139] en_b 
+ precharge 
* No parameters

xprecharge_140 
+ vdd bl[140] br[140] en_b 
+ precharge 
* No parameters

xprecharge_141 
+ vdd bl[141] br[141] en_b 
+ precharge 
* No parameters

xprecharge_142 
+ vdd bl[142] br[142] en_b 
+ precharge 
* No parameters

xprecharge_143 
+ vdd bl[143] br[143] en_b 
+ precharge 
* No parameters

xprecharge_144 
+ vdd bl[144] br[144] en_b 
+ precharge 
* No parameters

xprecharge_145 
+ vdd bl[145] br[145] en_b 
+ precharge 
* No parameters

xprecharge_146 
+ vdd bl[146] br[146] en_b 
+ precharge 
* No parameters

xprecharge_147 
+ vdd bl[147] br[147] en_b 
+ precharge 
* No parameters

xprecharge_148 
+ vdd bl[148] br[148] en_b 
+ precharge 
* No parameters

xprecharge_149 
+ vdd bl[149] br[149] en_b 
+ precharge 
* No parameters

xprecharge_150 
+ vdd bl[150] br[150] en_b 
+ precharge 
* No parameters

xprecharge_151 
+ vdd bl[151] br[151] en_b 
+ precharge 
* No parameters

xprecharge_152 
+ vdd bl[152] br[152] en_b 
+ precharge 
* No parameters

xprecharge_153 
+ vdd bl[153] br[153] en_b 
+ precharge 
* No parameters

xprecharge_154 
+ vdd bl[154] br[154] en_b 
+ precharge 
* No parameters

xprecharge_155 
+ vdd bl[155] br[155] en_b 
+ precharge 
* No parameters

xprecharge_156 
+ vdd bl[156] br[156] en_b 
+ precharge 
* No parameters

xprecharge_157 
+ vdd bl[157] br[157] en_b 
+ precharge 
* No parameters

xprecharge_158 
+ vdd bl[158] br[158] en_b 
+ precharge 
* No parameters

xprecharge_159 
+ vdd bl[159] br[159] en_b 
+ precharge 
* No parameters

xprecharge_160 
+ vdd bl[160] br[160] en_b 
+ precharge 
* No parameters

xprecharge_161 
+ vdd bl[161] br[161] en_b 
+ precharge 
* No parameters

xprecharge_162 
+ vdd bl[162] br[162] en_b 
+ precharge 
* No parameters

xprecharge_163 
+ vdd bl[163] br[163] en_b 
+ precharge 
* No parameters

xprecharge_164 
+ vdd bl[164] br[164] en_b 
+ precharge 
* No parameters

xprecharge_165 
+ vdd bl[165] br[165] en_b 
+ precharge 
* No parameters

xprecharge_166 
+ vdd bl[166] br[166] en_b 
+ precharge 
* No parameters

xprecharge_167 
+ vdd bl[167] br[167] en_b 
+ precharge 
* No parameters

xprecharge_168 
+ vdd bl[168] br[168] en_b 
+ precharge 
* No parameters

xprecharge_169 
+ vdd bl[169] br[169] en_b 
+ precharge 
* No parameters

xprecharge_170 
+ vdd bl[170] br[170] en_b 
+ precharge 
* No parameters

xprecharge_171 
+ vdd bl[171] br[171] en_b 
+ precharge 
* No parameters

xprecharge_172 
+ vdd bl[172] br[172] en_b 
+ precharge 
* No parameters

xprecharge_173 
+ vdd bl[173] br[173] en_b 
+ precharge 
* No parameters

xprecharge_174 
+ vdd bl[174] br[174] en_b 
+ precharge 
* No parameters

xprecharge_175 
+ vdd bl[175] br[175] en_b 
+ precharge 
* No parameters

xprecharge_176 
+ vdd bl[176] br[176] en_b 
+ precharge 
* No parameters

xprecharge_177 
+ vdd bl[177] br[177] en_b 
+ precharge 
* No parameters

xprecharge_178 
+ vdd bl[178] br[178] en_b 
+ precharge 
* No parameters

xprecharge_179 
+ vdd bl[179] br[179] en_b 
+ precharge 
* No parameters

xprecharge_180 
+ vdd bl[180] br[180] en_b 
+ precharge 
* No parameters

xprecharge_181 
+ vdd bl[181] br[181] en_b 
+ precharge 
* No parameters

xprecharge_182 
+ vdd bl[182] br[182] en_b 
+ precharge 
* No parameters

xprecharge_183 
+ vdd bl[183] br[183] en_b 
+ precharge 
* No parameters

xprecharge_184 
+ vdd bl[184] br[184] en_b 
+ precharge 
* No parameters

xprecharge_185 
+ vdd bl[185] br[185] en_b 
+ precharge 
* No parameters

xprecharge_186 
+ vdd bl[186] br[186] en_b 
+ precharge 
* No parameters

xprecharge_187 
+ vdd bl[187] br[187] en_b 
+ precharge 
* No parameters

xprecharge_188 
+ vdd bl[188] br[188] en_b 
+ precharge 
* No parameters

xprecharge_189 
+ vdd bl[189] br[189] en_b 
+ precharge 
* No parameters

xprecharge_190 
+ vdd bl[190] br[190] en_b 
+ precharge 
* No parameters

xprecharge_191 
+ vdd bl[191] br[191] en_b 
+ precharge 
* No parameters

xprecharge_192 
+ vdd bl[192] br[192] en_b 
+ precharge 
* No parameters

xprecharge_193 
+ vdd bl[193] br[193] en_b 
+ precharge 
* No parameters

xprecharge_194 
+ vdd bl[194] br[194] en_b 
+ precharge 
* No parameters

xprecharge_195 
+ vdd bl[195] br[195] en_b 
+ precharge 
* No parameters

xprecharge_196 
+ vdd bl[196] br[196] en_b 
+ precharge 
* No parameters

xprecharge_197 
+ vdd bl[197] br[197] en_b 
+ precharge 
* No parameters

xprecharge_198 
+ vdd bl[198] br[198] en_b 
+ precharge 
* No parameters

xprecharge_199 
+ vdd bl[199] br[199] en_b 
+ precharge 
* No parameters

xprecharge_200 
+ vdd bl[200] br[200] en_b 
+ precharge 
* No parameters

xprecharge_201 
+ vdd bl[201] br[201] en_b 
+ precharge 
* No parameters

xprecharge_202 
+ vdd bl[202] br[202] en_b 
+ precharge 
* No parameters

xprecharge_203 
+ vdd bl[203] br[203] en_b 
+ precharge 
* No parameters

xprecharge_204 
+ vdd bl[204] br[204] en_b 
+ precharge 
* No parameters

xprecharge_205 
+ vdd bl[205] br[205] en_b 
+ precharge 
* No parameters

xprecharge_206 
+ vdd bl[206] br[206] en_b 
+ precharge 
* No parameters

xprecharge_207 
+ vdd bl[207] br[207] en_b 
+ precharge 
* No parameters

xprecharge_208 
+ vdd bl[208] br[208] en_b 
+ precharge 
* No parameters

xprecharge_209 
+ vdd bl[209] br[209] en_b 
+ precharge 
* No parameters

xprecharge_210 
+ vdd bl[210] br[210] en_b 
+ precharge 
* No parameters

xprecharge_211 
+ vdd bl[211] br[211] en_b 
+ precharge 
* No parameters

xprecharge_212 
+ vdd bl[212] br[212] en_b 
+ precharge 
* No parameters

xprecharge_213 
+ vdd bl[213] br[213] en_b 
+ precharge 
* No parameters

xprecharge_214 
+ vdd bl[214] br[214] en_b 
+ precharge 
* No parameters

xprecharge_215 
+ vdd bl[215] br[215] en_b 
+ precharge 
* No parameters

xprecharge_216 
+ vdd bl[216] br[216] en_b 
+ precharge 
* No parameters

xprecharge_217 
+ vdd bl[217] br[217] en_b 
+ precharge 
* No parameters

xprecharge_218 
+ vdd bl[218] br[218] en_b 
+ precharge 
* No parameters

xprecharge_219 
+ vdd bl[219] br[219] en_b 
+ precharge 
* No parameters

xprecharge_220 
+ vdd bl[220] br[220] en_b 
+ precharge 
* No parameters

xprecharge_221 
+ vdd bl[221] br[221] en_b 
+ precharge 
* No parameters

xprecharge_222 
+ vdd bl[222] br[222] en_b 
+ precharge 
* No parameters

xprecharge_223 
+ vdd bl[223] br[223] en_b 
+ precharge 
* No parameters

xprecharge_224 
+ vdd bl[224] br[224] en_b 
+ precharge 
* No parameters

xprecharge_225 
+ vdd bl[225] br[225] en_b 
+ precharge 
* No parameters

xprecharge_226 
+ vdd bl[226] br[226] en_b 
+ precharge 
* No parameters

xprecharge_227 
+ vdd bl[227] br[227] en_b 
+ precharge 
* No parameters

xprecharge_228 
+ vdd bl[228] br[228] en_b 
+ precharge 
* No parameters

xprecharge_229 
+ vdd bl[229] br[229] en_b 
+ precharge 
* No parameters

xprecharge_230 
+ vdd bl[230] br[230] en_b 
+ precharge 
* No parameters

xprecharge_231 
+ vdd bl[231] br[231] en_b 
+ precharge 
* No parameters

xprecharge_232 
+ vdd bl[232] br[232] en_b 
+ precharge 
* No parameters

xprecharge_233 
+ vdd bl[233] br[233] en_b 
+ precharge 
* No parameters

xprecharge_234 
+ vdd bl[234] br[234] en_b 
+ precharge 
* No parameters

xprecharge_235 
+ vdd bl[235] br[235] en_b 
+ precharge 
* No parameters

xprecharge_236 
+ vdd bl[236] br[236] en_b 
+ precharge 
* No parameters

xprecharge_237 
+ vdd bl[237] br[237] en_b 
+ precharge 
* No parameters

xprecharge_238 
+ vdd bl[238] br[238] en_b 
+ precharge 
* No parameters

xprecharge_239 
+ vdd bl[239] br[239] en_b 
+ precharge 
* No parameters

xprecharge_240 
+ vdd bl[240] br[240] en_b 
+ precharge 
* No parameters

xprecharge_241 
+ vdd bl[241] br[241] en_b 
+ precharge 
* No parameters

xprecharge_242 
+ vdd bl[242] br[242] en_b 
+ precharge 
* No parameters

xprecharge_243 
+ vdd bl[243] br[243] en_b 
+ precharge 
* No parameters

xprecharge_244 
+ vdd bl[244] br[244] en_b 
+ precharge 
* No parameters

xprecharge_245 
+ vdd bl[245] br[245] en_b 
+ precharge 
* No parameters

xprecharge_246 
+ vdd bl[246] br[246] en_b 
+ precharge 
* No parameters

xprecharge_247 
+ vdd bl[247] br[247] en_b 
+ precharge 
* No parameters

xprecharge_248 
+ vdd bl[248] br[248] en_b 
+ precharge 
* No parameters

xprecharge_249 
+ vdd bl[249] br[249] en_b 
+ precharge 
* No parameters

xprecharge_250 
+ vdd bl[250] br[250] en_b 
+ precharge 
* No parameters

xprecharge_251 
+ vdd bl[251] br[251] en_b 
+ precharge 
* No parameters

xprecharge_252 
+ vdd bl[252] br[252] en_b 
+ precharge 
* No parameters

xprecharge_253 
+ vdd bl[253] br[253] en_b 
+ precharge 
* No parameters

xprecharge_254 
+ vdd bl[254] br[254] en_b 
+ precharge 
* No parameters

xprecharge_255 
+ vdd bl[255] br[255] en_b 
+ precharge 
* No parameters

xprecharge_256 
+ vdd bl[256] br[256] en_b 
+ precharge 
* No parameters

.ENDS

.SUBCKT read_mux 
+ sel_b bl br bl_out br_out vdd 

xMBL 
+ bl_out sel_b bl vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

xMBR 
+ br_out sel_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

.ENDS

.SUBCKT read_mux_array 
+ sel_b[7] sel_b[6] sel_b[5] sel_b[4] sel_b[3] sel_b[2] sel_b[1] sel_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_out[31] bl_out[30] bl_out[29] bl_out[28] bl_out[27] bl_out[26] bl_out[25] bl_out[24] bl_out[23] bl_out[22] bl_out[21] bl_out[20] bl_out[19] bl_out[18] bl_out[17] bl_out[16] bl_out[15] bl_out[14] bl_out[13] bl_out[12] bl_out[11] bl_out[10] bl_out[9] bl_out[8] bl_out[7] bl_out[6] bl_out[5] bl_out[4] bl_out[3] bl_out[2] bl_out[1] bl_out[0] br_out[31] br_out[30] br_out[29] br_out[28] br_out[27] br_out[26] br_out[25] br_out[24] br_out[23] br_out[22] br_out[21] br_out[20] br_out[19] br_out[18] br_out[17] br_out[16] br_out[15] br_out[14] br_out[13] br_out[12] br_out[11] br_out[10] br_out[9] br_out[8] br_out[7] br_out[6] br_out[5] br_out[4] br_out[3] br_out[2] br_out[1] br_out[0] vdd 

xmux_0 
+ sel_b[0] bl[0] br[0] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_1 
+ sel_b[1] bl[1] br[1] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_2 
+ sel_b[2] bl[2] br[2] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_3 
+ sel_b[3] bl[3] br[3] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_4 
+ sel_b[4] bl[4] br[4] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_5 
+ sel_b[5] bl[5] br[5] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_6 
+ sel_b[6] bl[6] br[6] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_7 
+ sel_b[7] bl[7] br[7] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_8 
+ sel_b[0] bl[8] br[8] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_9 
+ sel_b[1] bl[9] br[9] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_10 
+ sel_b[2] bl[10] br[10] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_11 
+ sel_b[3] bl[11] br[11] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_12 
+ sel_b[4] bl[12] br[12] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_13 
+ sel_b[5] bl[13] br[13] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_14 
+ sel_b[6] bl[14] br[14] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_15 
+ sel_b[7] bl[15] br[15] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_16 
+ sel_b[0] bl[16] br[16] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_17 
+ sel_b[1] bl[17] br[17] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_18 
+ sel_b[2] bl[18] br[18] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_19 
+ sel_b[3] bl[19] br[19] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_20 
+ sel_b[4] bl[20] br[20] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_21 
+ sel_b[5] bl[21] br[21] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_22 
+ sel_b[6] bl[22] br[22] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_23 
+ sel_b[7] bl[23] br[23] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_24 
+ sel_b[0] bl[24] br[24] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_25 
+ sel_b[1] bl[25] br[25] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_26 
+ sel_b[2] bl[26] br[26] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_27 
+ sel_b[3] bl[27] br[27] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_28 
+ sel_b[4] bl[28] br[28] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_29 
+ sel_b[5] bl[29] br[29] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_30 
+ sel_b[6] bl[30] br[30] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_31 
+ sel_b[7] bl[31] br[31] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_32 
+ sel_b[0] bl[32] br[32] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_33 
+ sel_b[1] bl[33] br[33] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_34 
+ sel_b[2] bl[34] br[34] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_35 
+ sel_b[3] bl[35] br[35] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_36 
+ sel_b[4] bl[36] br[36] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_37 
+ sel_b[5] bl[37] br[37] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_38 
+ sel_b[6] bl[38] br[38] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_39 
+ sel_b[7] bl[39] br[39] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_40 
+ sel_b[0] bl[40] br[40] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_41 
+ sel_b[1] bl[41] br[41] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_42 
+ sel_b[2] bl[42] br[42] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_43 
+ sel_b[3] bl[43] br[43] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_44 
+ sel_b[4] bl[44] br[44] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_45 
+ sel_b[5] bl[45] br[45] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_46 
+ sel_b[6] bl[46] br[46] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_47 
+ sel_b[7] bl[47] br[47] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_48 
+ sel_b[0] bl[48] br[48] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_49 
+ sel_b[1] bl[49] br[49] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_50 
+ sel_b[2] bl[50] br[50] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_51 
+ sel_b[3] bl[51] br[51] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_52 
+ sel_b[4] bl[52] br[52] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_53 
+ sel_b[5] bl[53] br[53] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_54 
+ sel_b[6] bl[54] br[54] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_55 
+ sel_b[7] bl[55] br[55] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_56 
+ sel_b[0] bl[56] br[56] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_57 
+ sel_b[1] bl[57] br[57] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_58 
+ sel_b[2] bl[58] br[58] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_59 
+ sel_b[3] bl[59] br[59] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_60 
+ sel_b[4] bl[60] br[60] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_61 
+ sel_b[5] bl[61] br[61] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_62 
+ sel_b[6] bl[62] br[62] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_63 
+ sel_b[7] bl[63] br[63] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_64 
+ sel_b[0] bl[64] br[64] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_65 
+ sel_b[1] bl[65] br[65] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_66 
+ sel_b[2] bl[66] br[66] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_67 
+ sel_b[3] bl[67] br[67] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_68 
+ sel_b[4] bl[68] br[68] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_69 
+ sel_b[5] bl[69] br[69] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_70 
+ sel_b[6] bl[70] br[70] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_71 
+ sel_b[7] bl[71] br[71] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_72 
+ sel_b[0] bl[72] br[72] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_73 
+ sel_b[1] bl[73] br[73] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_74 
+ sel_b[2] bl[74] br[74] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_75 
+ sel_b[3] bl[75] br[75] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_76 
+ sel_b[4] bl[76] br[76] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_77 
+ sel_b[5] bl[77] br[77] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_78 
+ sel_b[6] bl[78] br[78] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_79 
+ sel_b[7] bl[79] br[79] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_80 
+ sel_b[0] bl[80] br[80] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_81 
+ sel_b[1] bl[81] br[81] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_82 
+ sel_b[2] bl[82] br[82] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_83 
+ sel_b[3] bl[83] br[83] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_84 
+ sel_b[4] bl[84] br[84] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_85 
+ sel_b[5] bl[85] br[85] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_86 
+ sel_b[6] bl[86] br[86] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_87 
+ sel_b[7] bl[87] br[87] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_88 
+ sel_b[0] bl[88] br[88] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_89 
+ sel_b[1] bl[89] br[89] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_90 
+ sel_b[2] bl[90] br[90] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_91 
+ sel_b[3] bl[91] br[91] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_92 
+ sel_b[4] bl[92] br[92] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_93 
+ sel_b[5] bl[93] br[93] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_94 
+ sel_b[6] bl[94] br[94] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_95 
+ sel_b[7] bl[95] br[95] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_96 
+ sel_b[0] bl[96] br[96] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_97 
+ sel_b[1] bl[97] br[97] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_98 
+ sel_b[2] bl[98] br[98] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_99 
+ sel_b[3] bl[99] br[99] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_100 
+ sel_b[4] bl[100] br[100] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_101 
+ sel_b[5] bl[101] br[101] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_102 
+ sel_b[6] bl[102] br[102] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_103 
+ sel_b[7] bl[103] br[103] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_104 
+ sel_b[0] bl[104] br[104] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_105 
+ sel_b[1] bl[105] br[105] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_106 
+ sel_b[2] bl[106] br[106] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_107 
+ sel_b[3] bl[107] br[107] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_108 
+ sel_b[4] bl[108] br[108] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_109 
+ sel_b[5] bl[109] br[109] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_110 
+ sel_b[6] bl[110] br[110] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_111 
+ sel_b[7] bl[111] br[111] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_112 
+ sel_b[0] bl[112] br[112] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_113 
+ sel_b[1] bl[113] br[113] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_114 
+ sel_b[2] bl[114] br[114] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_115 
+ sel_b[3] bl[115] br[115] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_116 
+ sel_b[4] bl[116] br[116] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_117 
+ sel_b[5] bl[117] br[117] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_118 
+ sel_b[6] bl[118] br[118] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_119 
+ sel_b[7] bl[119] br[119] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_120 
+ sel_b[0] bl[120] br[120] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_121 
+ sel_b[1] bl[121] br[121] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_122 
+ sel_b[2] bl[122] br[122] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_123 
+ sel_b[3] bl[123] br[123] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_124 
+ sel_b[4] bl[124] br[124] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_125 
+ sel_b[5] bl[125] br[125] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_126 
+ sel_b[6] bl[126] br[126] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_127 
+ sel_b[7] bl[127] br[127] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_128 
+ sel_b[0] bl[128] br[128] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_129 
+ sel_b[1] bl[129] br[129] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_130 
+ sel_b[2] bl[130] br[130] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_131 
+ sel_b[3] bl[131] br[131] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_132 
+ sel_b[4] bl[132] br[132] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_133 
+ sel_b[5] bl[133] br[133] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_134 
+ sel_b[6] bl[134] br[134] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_135 
+ sel_b[7] bl[135] br[135] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_136 
+ sel_b[0] bl[136] br[136] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_137 
+ sel_b[1] bl[137] br[137] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_138 
+ sel_b[2] bl[138] br[138] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_139 
+ sel_b[3] bl[139] br[139] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_140 
+ sel_b[4] bl[140] br[140] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_141 
+ sel_b[5] bl[141] br[141] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_142 
+ sel_b[6] bl[142] br[142] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_143 
+ sel_b[7] bl[143] br[143] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_144 
+ sel_b[0] bl[144] br[144] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_145 
+ sel_b[1] bl[145] br[145] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_146 
+ sel_b[2] bl[146] br[146] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_147 
+ sel_b[3] bl[147] br[147] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_148 
+ sel_b[4] bl[148] br[148] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_149 
+ sel_b[5] bl[149] br[149] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_150 
+ sel_b[6] bl[150] br[150] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_151 
+ sel_b[7] bl[151] br[151] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_152 
+ sel_b[0] bl[152] br[152] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_153 
+ sel_b[1] bl[153] br[153] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_154 
+ sel_b[2] bl[154] br[154] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_155 
+ sel_b[3] bl[155] br[155] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_156 
+ sel_b[4] bl[156] br[156] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_157 
+ sel_b[5] bl[157] br[157] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_158 
+ sel_b[6] bl[158] br[158] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_159 
+ sel_b[7] bl[159] br[159] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_160 
+ sel_b[0] bl[160] br[160] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_161 
+ sel_b[1] bl[161] br[161] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_162 
+ sel_b[2] bl[162] br[162] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_163 
+ sel_b[3] bl[163] br[163] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_164 
+ sel_b[4] bl[164] br[164] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_165 
+ sel_b[5] bl[165] br[165] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_166 
+ sel_b[6] bl[166] br[166] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_167 
+ sel_b[7] bl[167] br[167] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_168 
+ sel_b[0] bl[168] br[168] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_169 
+ sel_b[1] bl[169] br[169] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_170 
+ sel_b[2] bl[170] br[170] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_171 
+ sel_b[3] bl[171] br[171] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_172 
+ sel_b[4] bl[172] br[172] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_173 
+ sel_b[5] bl[173] br[173] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_174 
+ sel_b[6] bl[174] br[174] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_175 
+ sel_b[7] bl[175] br[175] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_176 
+ sel_b[0] bl[176] br[176] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_177 
+ sel_b[1] bl[177] br[177] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_178 
+ sel_b[2] bl[178] br[178] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_179 
+ sel_b[3] bl[179] br[179] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_180 
+ sel_b[4] bl[180] br[180] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_181 
+ sel_b[5] bl[181] br[181] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_182 
+ sel_b[6] bl[182] br[182] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_183 
+ sel_b[7] bl[183] br[183] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_184 
+ sel_b[0] bl[184] br[184] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_185 
+ sel_b[1] bl[185] br[185] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_186 
+ sel_b[2] bl[186] br[186] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_187 
+ sel_b[3] bl[187] br[187] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_188 
+ sel_b[4] bl[188] br[188] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_189 
+ sel_b[5] bl[189] br[189] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_190 
+ sel_b[6] bl[190] br[190] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_191 
+ sel_b[7] bl[191] br[191] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_192 
+ sel_b[0] bl[192] br[192] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_193 
+ sel_b[1] bl[193] br[193] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_194 
+ sel_b[2] bl[194] br[194] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_195 
+ sel_b[3] bl[195] br[195] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_196 
+ sel_b[4] bl[196] br[196] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_197 
+ sel_b[5] bl[197] br[197] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_198 
+ sel_b[6] bl[198] br[198] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_199 
+ sel_b[7] bl[199] br[199] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_200 
+ sel_b[0] bl[200] br[200] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_201 
+ sel_b[1] bl[201] br[201] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_202 
+ sel_b[2] bl[202] br[202] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_203 
+ sel_b[3] bl[203] br[203] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_204 
+ sel_b[4] bl[204] br[204] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_205 
+ sel_b[5] bl[205] br[205] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_206 
+ sel_b[6] bl[206] br[206] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_207 
+ sel_b[7] bl[207] br[207] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_208 
+ sel_b[0] bl[208] br[208] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_209 
+ sel_b[1] bl[209] br[209] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_210 
+ sel_b[2] bl[210] br[210] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_211 
+ sel_b[3] bl[211] br[211] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_212 
+ sel_b[4] bl[212] br[212] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_213 
+ sel_b[5] bl[213] br[213] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_214 
+ sel_b[6] bl[214] br[214] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_215 
+ sel_b[7] bl[215] br[215] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_216 
+ sel_b[0] bl[216] br[216] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_217 
+ sel_b[1] bl[217] br[217] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_218 
+ sel_b[2] bl[218] br[218] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_219 
+ sel_b[3] bl[219] br[219] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_220 
+ sel_b[4] bl[220] br[220] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_221 
+ sel_b[5] bl[221] br[221] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_222 
+ sel_b[6] bl[222] br[222] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_223 
+ sel_b[7] bl[223] br[223] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_224 
+ sel_b[0] bl[224] br[224] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_225 
+ sel_b[1] bl[225] br[225] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_226 
+ sel_b[2] bl[226] br[226] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_227 
+ sel_b[3] bl[227] br[227] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_228 
+ sel_b[4] bl[228] br[228] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_229 
+ sel_b[5] bl[229] br[229] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_230 
+ sel_b[6] bl[230] br[230] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_231 
+ sel_b[7] bl[231] br[231] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_232 
+ sel_b[0] bl[232] br[232] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_233 
+ sel_b[1] bl[233] br[233] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_234 
+ sel_b[2] bl[234] br[234] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_235 
+ sel_b[3] bl[235] br[235] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_236 
+ sel_b[4] bl[236] br[236] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_237 
+ sel_b[5] bl[237] br[237] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_238 
+ sel_b[6] bl[238] br[238] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_239 
+ sel_b[7] bl[239] br[239] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_240 
+ sel_b[0] bl[240] br[240] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_241 
+ sel_b[1] bl[241] br[241] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_242 
+ sel_b[2] bl[242] br[242] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_243 
+ sel_b[3] bl[243] br[243] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_244 
+ sel_b[4] bl[244] br[244] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_245 
+ sel_b[5] bl[245] br[245] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_246 
+ sel_b[6] bl[246] br[246] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_247 
+ sel_b[7] bl[247] br[247] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_248 
+ sel_b[0] bl[248] br[248] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_249 
+ sel_b[1] bl[249] br[249] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_250 
+ sel_b[2] bl[250] br[250] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_251 
+ sel_b[3] bl[251] br[251] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_252 
+ sel_b[4] bl[252] br[252] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_253 
+ sel_b[5] bl[253] br[253] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_254 
+ sel_b[6] bl[254] br[254] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_255 
+ sel_b[7] bl[255] br[255] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

.ENDS

.SUBCKT write_mux 
+ we data data_b bl br vss 

xMMUXBR 
+ br data x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMMUXBL 
+ bl data_b x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMPD 
+ x we vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT write_mux_array 
+ we[7] we[6] we[5] we[4] we[3] we[2] we[1] we[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 

xmux_0 
+ we[0] data[0] data_b[0] bl[0] br[0] vss 
+ write_mux 
* No parameters

xmux_1 
+ we[1] data[0] data_b[0] bl[1] br[1] vss 
+ write_mux 
* No parameters

xmux_2 
+ we[2] data[0] data_b[0] bl[2] br[2] vss 
+ write_mux 
* No parameters

xmux_3 
+ we[3] data[0] data_b[0] bl[3] br[3] vss 
+ write_mux 
* No parameters

xmux_4 
+ we[4] data[0] data_b[0] bl[4] br[4] vss 
+ write_mux 
* No parameters

xmux_5 
+ we[5] data[0] data_b[0] bl[5] br[5] vss 
+ write_mux 
* No parameters

xmux_6 
+ we[6] data[0] data_b[0] bl[6] br[6] vss 
+ write_mux 
* No parameters

xmux_7 
+ we[7] data[0] data_b[0] bl[7] br[7] vss 
+ write_mux 
* No parameters

xmux_8 
+ we[0] data[1] data_b[1] bl[8] br[8] vss 
+ write_mux 
* No parameters

xmux_9 
+ we[1] data[1] data_b[1] bl[9] br[9] vss 
+ write_mux 
* No parameters

xmux_10 
+ we[2] data[1] data_b[1] bl[10] br[10] vss 
+ write_mux 
* No parameters

xmux_11 
+ we[3] data[1] data_b[1] bl[11] br[11] vss 
+ write_mux 
* No parameters

xmux_12 
+ we[4] data[1] data_b[1] bl[12] br[12] vss 
+ write_mux 
* No parameters

xmux_13 
+ we[5] data[1] data_b[1] bl[13] br[13] vss 
+ write_mux 
* No parameters

xmux_14 
+ we[6] data[1] data_b[1] bl[14] br[14] vss 
+ write_mux 
* No parameters

xmux_15 
+ we[7] data[1] data_b[1] bl[15] br[15] vss 
+ write_mux 
* No parameters

xmux_16 
+ we[0] data[2] data_b[2] bl[16] br[16] vss 
+ write_mux 
* No parameters

xmux_17 
+ we[1] data[2] data_b[2] bl[17] br[17] vss 
+ write_mux 
* No parameters

xmux_18 
+ we[2] data[2] data_b[2] bl[18] br[18] vss 
+ write_mux 
* No parameters

xmux_19 
+ we[3] data[2] data_b[2] bl[19] br[19] vss 
+ write_mux 
* No parameters

xmux_20 
+ we[4] data[2] data_b[2] bl[20] br[20] vss 
+ write_mux 
* No parameters

xmux_21 
+ we[5] data[2] data_b[2] bl[21] br[21] vss 
+ write_mux 
* No parameters

xmux_22 
+ we[6] data[2] data_b[2] bl[22] br[22] vss 
+ write_mux 
* No parameters

xmux_23 
+ we[7] data[2] data_b[2] bl[23] br[23] vss 
+ write_mux 
* No parameters

xmux_24 
+ we[0] data[3] data_b[3] bl[24] br[24] vss 
+ write_mux 
* No parameters

xmux_25 
+ we[1] data[3] data_b[3] bl[25] br[25] vss 
+ write_mux 
* No parameters

xmux_26 
+ we[2] data[3] data_b[3] bl[26] br[26] vss 
+ write_mux 
* No parameters

xmux_27 
+ we[3] data[3] data_b[3] bl[27] br[27] vss 
+ write_mux 
* No parameters

xmux_28 
+ we[4] data[3] data_b[3] bl[28] br[28] vss 
+ write_mux 
* No parameters

xmux_29 
+ we[5] data[3] data_b[3] bl[29] br[29] vss 
+ write_mux 
* No parameters

xmux_30 
+ we[6] data[3] data_b[3] bl[30] br[30] vss 
+ write_mux 
* No parameters

xmux_31 
+ we[7] data[3] data_b[3] bl[31] br[31] vss 
+ write_mux 
* No parameters

xmux_32 
+ we[0] data[4] data_b[4] bl[32] br[32] vss 
+ write_mux 
* No parameters

xmux_33 
+ we[1] data[4] data_b[4] bl[33] br[33] vss 
+ write_mux 
* No parameters

xmux_34 
+ we[2] data[4] data_b[4] bl[34] br[34] vss 
+ write_mux 
* No parameters

xmux_35 
+ we[3] data[4] data_b[4] bl[35] br[35] vss 
+ write_mux 
* No parameters

xmux_36 
+ we[4] data[4] data_b[4] bl[36] br[36] vss 
+ write_mux 
* No parameters

xmux_37 
+ we[5] data[4] data_b[4] bl[37] br[37] vss 
+ write_mux 
* No parameters

xmux_38 
+ we[6] data[4] data_b[4] bl[38] br[38] vss 
+ write_mux 
* No parameters

xmux_39 
+ we[7] data[4] data_b[4] bl[39] br[39] vss 
+ write_mux 
* No parameters

xmux_40 
+ we[0] data[5] data_b[5] bl[40] br[40] vss 
+ write_mux 
* No parameters

xmux_41 
+ we[1] data[5] data_b[5] bl[41] br[41] vss 
+ write_mux 
* No parameters

xmux_42 
+ we[2] data[5] data_b[5] bl[42] br[42] vss 
+ write_mux 
* No parameters

xmux_43 
+ we[3] data[5] data_b[5] bl[43] br[43] vss 
+ write_mux 
* No parameters

xmux_44 
+ we[4] data[5] data_b[5] bl[44] br[44] vss 
+ write_mux 
* No parameters

xmux_45 
+ we[5] data[5] data_b[5] bl[45] br[45] vss 
+ write_mux 
* No parameters

xmux_46 
+ we[6] data[5] data_b[5] bl[46] br[46] vss 
+ write_mux 
* No parameters

xmux_47 
+ we[7] data[5] data_b[5] bl[47] br[47] vss 
+ write_mux 
* No parameters

xmux_48 
+ we[0] data[6] data_b[6] bl[48] br[48] vss 
+ write_mux 
* No parameters

xmux_49 
+ we[1] data[6] data_b[6] bl[49] br[49] vss 
+ write_mux 
* No parameters

xmux_50 
+ we[2] data[6] data_b[6] bl[50] br[50] vss 
+ write_mux 
* No parameters

xmux_51 
+ we[3] data[6] data_b[6] bl[51] br[51] vss 
+ write_mux 
* No parameters

xmux_52 
+ we[4] data[6] data_b[6] bl[52] br[52] vss 
+ write_mux 
* No parameters

xmux_53 
+ we[5] data[6] data_b[6] bl[53] br[53] vss 
+ write_mux 
* No parameters

xmux_54 
+ we[6] data[6] data_b[6] bl[54] br[54] vss 
+ write_mux 
* No parameters

xmux_55 
+ we[7] data[6] data_b[6] bl[55] br[55] vss 
+ write_mux 
* No parameters

xmux_56 
+ we[0] data[7] data_b[7] bl[56] br[56] vss 
+ write_mux 
* No parameters

xmux_57 
+ we[1] data[7] data_b[7] bl[57] br[57] vss 
+ write_mux 
* No parameters

xmux_58 
+ we[2] data[7] data_b[7] bl[58] br[58] vss 
+ write_mux 
* No parameters

xmux_59 
+ we[3] data[7] data_b[7] bl[59] br[59] vss 
+ write_mux 
* No parameters

xmux_60 
+ we[4] data[7] data_b[7] bl[60] br[60] vss 
+ write_mux 
* No parameters

xmux_61 
+ we[5] data[7] data_b[7] bl[61] br[61] vss 
+ write_mux 
* No parameters

xmux_62 
+ we[6] data[7] data_b[7] bl[62] br[62] vss 
+ write_mux 
* No parameters

xmux_63 
+ we[7] data[7] data_b[7] bl[63] br[63] vss 
+ write_mux 
* No parameters

xmux_64 
+ we[0] data[8] data_b[8] bl[64] br[64] vss 
+ write_mux 
* No parameters

xmux_65 
+ we[1] data[8] data_b[8] bl[65] br[65] vss 
+ write_mux 
* No parameters

xmux_66 
+ we[2] data[8] data_b[8] bl[66] br[66] vss 
+ write_mux 
* No parameters

xmux_67 
+ we[3] data[8] data_b[8] bl[67] br[67] vss 
+ write_mux 
* No parameters

xmux_68 
+ we[4] data[8] data_b[8] bl[68] br[68] vss 
+ write_mux 
* No parameters

xmux_69 
+ we[5] data[8] data_b[8] bl[69] br[69] vss 
+ write_mux 
* No parameters

xmux_70 
+ we[6] data[8] data_b[8] bl[70] br[70] vss 
+ write_mux 
* No parameters

xmux_71 
+ we[7] data[8] data_b[8] bl[71] br[71] vss 
+ write_mux 
* No parameters

xmux_72 
+ we[0] data[9] data_b[9] bl[72] br[72] vss 
+ write_mux 
* No parameters

xmux_73 
+ we[1] data[9] data_b[9] bl[73] br[73] vss 
+ write_mux 
* No parameters

xmux_74 
+ we[2] data[9] data_b[9] bl[74] br[74] vss 
+ write_mux 
* No parameters

xmux_75 
+ we[3] data[9] data_b[9] bl[75] br[75] vss 
+ write_mux 
* No parameters

xmux_76 
+ we[4] data[9] data_b[9] bl[76] br[76] vss 
+ write_mux 
* No parameters

xmux_77 
+ we[5] data[9] data_b[9] bl[77] br[77] vss 
+ write_mux 
* No parameters

xmux_78 
+ we[6] data[9] data_b[9] bl[78] br[78] vss 
+ write_mux 
* No parameters

xmux_79 
+ we[7] data[9] data_b[9] bl[79] br[79] vss 
+ write_mux 
* No parameters

xmux_80 
+ we[0] data[10] data_b[10] bl[80] br[80] vss 
+ write_mux 
* No parameters

xmux_81 
+ we[1] data[10] data_b[10] bl[81] br[81] vss 
+ write_mux 
* No parameters

xmux_82 
+ we[2] data[10] data_b[10] bl[82] br[82] vss 
+ write_mux 
* No parameters

xmux_83 
+ we[3] data[10] data_b[10] bl[83] br[83] vss 
+ write_mux 
* No parameters

xmux_84 
+ we[4] data[10] data_b[10] bl[84] br[84] vss 
+ write_mux 
* No parameters

xmux_85 
+ we[5] data[10] data_b[10] bl[85] br[85] vss 
+ write_mux 
* No parameters

xmux_86 
+ we[6] data[10] data_b[10] bl[86] br[86] vss 
+ write_mux 
* No parameters

xmux_87 
+ we[7] data[10] data_b[10] bl[87] br[87] vss 
+ write_mux 
* No parameters

xmux_88 
+ we[0] data[11] data_b[11] bl[88] br[88] vss 
+ write_mux 
* No parameters

xmux_89 
+ we[1] data[11] data_b[11] bl[89] br[89] vss 
+ write_mux 
* No parameters

xmux_90 
+ we[2] data[11] data_b[11] bl[90] br[90] vss 
+ write_mux 
* No parameters

xmux_91 
+ we[3] data[11] data_b[11] bl[91] br[91] vss 
+ write_mux 
* No parameters

xmux_92 
+ we[4] data[11] data_b[11] bl[92] br[92] vss 
+ write_mux 
* No parameters

xmux_93 
+ we[5] data[11] data_b[11] bl[93] br[93] vss 
+ write_mux 
* No parameters

xmux_94 
+ we[6] data[11] data_b[11] bl[94] br[94] vss 
+ write_mux 
* No parameters

xmux_95 
+ we[7] data[11] data_b[11] bl[95] br[95] vss 
+ write_mux 
* No parameters

xmux_96 
+ we[0] data[12] data_b[12] bl[96] br[96] vss 
+ write_mux 
* No parameters

xmux_97 
+ we[1] data[12] data_b[12] bl[97] br[97] vss 
+ write_mux 
* No parameters

xmux_98 
+ we[2] data[12] data_b[12] bl[98] br[98] vss 
+ write_mux 
* No parameters

xmux_99 
+ we[3] data[12] data_b[12] bl[99] br[99] vss 
+ write_mux 
* No parameters

xmux_100 
+ we[4] data[12] data_b[12] bl[100] br[100] vss 
+ write_mux 
* No parameters

xmux_101 
+ we[5] data[12] data_b[12] bl[101] br[101] vss 
+ write_mux 
* No parameters

xmux_102 
+ we[6] data[12] data_b[12] bl[102] br[102] vss 
+ write_mux 
* No parameters

xmux_103 
+ we[7] data[12] data_b[12] bl[103] br[103] vss 
+ write_mux 
* No parameters

xmux_104 
+ we[0] data[13] data_b[13] bl[104] br[104] vss 
+ write_mux 
* No parameters

xmux_105 
+ we[1] data[13] data_b[13] bl[105] br[105] vss 
+ write_mux 
* No parameters

xmux_106 
+ we[2] data[13] data_b[13] bl[106] br[106] vss 
+ write_mux 
* No parameters

xmux_107 
+ we[3] data[13] data_b[13] bl[107] br[107] vss 
+ write_mux 
* No parameters

xmux_108 
+ we[4] data[13] data_b[13] bl[108] br[108] vss 
+ write_mux 
* No parameters

xmux_109 
+ we[5] data[13] data_b[13] bl[109] br[109] vss 
+ write_mux 
* No parameters

xmux_110 
+ we[6] data[13] data_b[13] bl[110] br[110] vss 
+ write_mux 
* No parameters

xmux_111 
+ we[7] data[13] data_b[13] bl[111] br[111] vss 
+ write_mux 
* No parameters

xmux_112 
+ we[0] data[14] data_b[14] bl[112] br[112] vss 
+ write_mux 
* No parameters

xmux_113 
+ we[1] data[14] data_b[14] bl[113] br[113] vss 
+ write_mux 
* No parameters

xmux_114 
+ we[2] data[14] data_b[14] bl[114] br[114] vss 
+ write_mux 
* No parameters

xmux_115 
+ we[3] data[14] data_b[14] bl[115] br[115] vss 
+ write_mux 
* No parameters

xmux_116 
+ we[4] data[14] data_b[14] bl[116] br[116] vss 
+ write_mux 
* No parameters

xmux_117 
+ we[5] data[14] data_b[14] bl[117] br[117] vss 
+ write_mux 
* No parameters

xmux_118 
+ we[6] data[14] data_b[14] bl[118] br[118] vss 
+ write_mux 
* No parameters

xmux_119 
+ we[7] data[14] data_b[14] bl[119] br[119] vss 
+ write_mux 
* No parameters

xmux_120 
+ we[0] data[15] data_b[15] bl[120] br[120] vss 
+ write_mux 
* No parameters

xmux_121 
+ we[1] data[15] data_b[15] bl[121] br[121] vss 
+ write_mux 
* No parameters

xmux_122 
+ we[2] data[15] data_b[15] bl[122] br[122] vss 
+ write_mux 
* No parameters

xmux_123 
+ we[3] data[15] data_b[15] bl[123] br[123] vss 
+ write_mux 
* No parameters

xmux_124 
+ we[4] data[15] data_b[15] bl[124] br[124] vss 
+ write_mux 
* No parameters

xmux_125 
+ we[5] data[15] data_b[15] bl[125] br[125] vss 
+ write_mux 
* No parameters

xmux_126 
+ we[6] data[15] data_b[15] bl[126] br[126] vss 
+ write_mux 
* No parameters

xmux_127 
+ we[7] data[15] data_b[15] bl[127] br[127] vss 
+ write_mux 
* No parameters

xmux_128 
+ we[0] data[16] data_b[16] bl[128] br[128] vss 
+ write_mux 
* No parameters

xmux_129 
+ we[1] data[16] data_b[16] bl[129] br[129] vss 
+ write_mux 
* No parameters

xmux_130 
+ we[2] data[16] data_b[16] bl[130] br[130] vss 
+ write_mux 
* No parameters

xmux_131 
+ we[3] data[16] data_b[16] bl[131] br[131] vss 
+ write_mux 
* No parameters

xmux_132 
+ we[4] data[16] data_b[16] bl[132] br[132] vss 
+ write_mux 
* No parameters

xmux_133 
+ we[5] data[16] data_b[16] bl[133] br[133] vss 
+ write_mux 
* No parameters

xmux_134 
+ we[6] data[16] data_b[16] bl[134] br[134] vss 
+ write_mux 
* No parameters

xmux_135 
+ we[7] data[16] data_b[16] bl[135] br[135] vss 
+ write_mux 
* No parameters

xmux_136 
+ we[0] data[17] data_b[17] bl[136] br[136] vss 
+ write_mux 
* No parameters

xmux_137 
+ we[1] data[17] data_b[17] bl[137] br[137] vss 
+ write_mux 
* No parameters

xmux_138 
+ we[2] data[17] data_b[17] bl[138] br[138] vss 
+ write_mux 
* No parameters

xmux_139 
+ we[3] data[17] data_b[17] bl[139] br[139] vss 
+ write_mux 
* No parameters

xmux_140 
+ we[4] data[17] data_b[17] bl[140] br[140] vss 
+ write_mux 
* No parameters

xmux_141 
+ we[5] data[17] data_b[17] bl[141] br[141] vss 
+ write_mux 
* No parameters

xmux_142 
+ we[6] data[17] data_b[17] bl[142] br[142] vss 
+ write_mux 
* No parameters

xmux_143 
+ we[7] data[17] data_b[17] bl[143] br[143] vss 
+ write_mux 
* No parameters

xmux_144 
+ we[0] data[18] data_b[18] bl[144] br[144] vss 
+ write_mux 
* No parameters

xmux_145 
+ we[1] data[18] data_b[18] bl[145] br[145] vss 
+ write_mux 
* No parameters

xmux_146 
+ we[2] data[18] data_b[18] bl[146] br[146] vss 
+ write_mux 
* No parameters

xmux_147 
+ we[3] data[18] data_b[18] bl[147] br[147] vss 
+ write_mux 
* No parameters

xmux_148 
+ we[4] data[18] data_b[18] bl[148] br[148] vss 
+ write_mux 
* No parameters

xmux_149 
+ we[5] data[18] data_b[18] bl[149] br[149] vss 
+ write_mux 
* No parameters

xmux_150 
+ we[6] data[18] data_b[18] bl[150] br[150] vss 
+ write_mux 
* No parameters

xmux_151 
+ we[7] data[18] data_b[18] bl[151] br[151] vss 
+ write_mux 
* No parameters

xmux_152 
+ we[0] data[19] data_b[19] bl[152] br[152] vss 
+ write_mux 
* No parameters

xmux_153 
+ we[1] data[19] data_b[19] bl[153] br[153] vss 
+ write_mux 
* No parameters

xmux_154 
+ we[2] data[19] data_b[19] bl[154] br[154] vss 
+ write_mux 
* No parameters

xmux_155 
+ we[3] data[19] data_b[19] bl[155] br[155] vss 
+ write_mux 
* No parameters

xmux_156 
+ we[4] data[19] data_b[19] bl[156] br[156] vss 
+ write_mux 
* No parameters

xmux_157 
+ we[5] data[19] data_b[19] bl[157] br[157] vss 
+ write_mux 
* No parameters

xmux_158 
+ we[6] data[19] data_b[19] bl[158] br[158] vss 
+ write_mux 
* No parameters

xmux_159 
+ we[7] data[19] data_b[19] bl[159] br[159] vss 
+ write_mux 
* No parameters

xmux_160 
+ we[0] data[20] data_b[20] bl[160] br[160] vss 
+ write_mux 
* No parameters

xmux_161 
+ we[1] data[20] data_b[20] bl[161] br[161] vss 
+ write_mux 
* No parameters

xmux_162 
+ we[2] data[20] data_b[20] bl[162] br[162] vss 
+ write_mux 
* No parameters

xmux_163 
+ we[3] data[20] data_b[20] bl[163] br[163] vss 
+ write_mux 
* No parameters

xmux_164 
+ we[4] data[20] data_b[20] bl[164] br[164] vss 
+ write_mux 
* No parameters

xmux_165 
+ we[5] data[20] data_b[20] bl[165] br[165] vss 
+ write_mux 
* No parameters

xmux_166 
+ we[6] data[20] data_b[20] bl[166] br[166] vss 
+ write_mux 
* No parameters

xmux_167 
+ we[7] data[20] data_b[20] bl[167] br[167] vss 
+ write_mux 
* No parameters

xmux_168 
+ we[0] data[21] data_b[21] bl[168] br[168] vss 
+ write_mux 
* No parameters

xmux_169 
+ we[1] data[21] data_b[21] bl[169] br[169] vss 
+ write_mux 
* No parameters

xmux_170 
+ we[2] data[21] data_b[21] bl[170] br[170] vss 
+ write_mux 
* No parameters

xmux_171 
+ we[3] data[21] data_b[21] bl[171] br[171] vss 
+ write_mux 
* No parameters

xmux_172 
+ we[4] data[21] data_b[21] bl[172] br[172] vss 
+ write_mux 
* No parameters

xmux_173 
+ we[5] data[21] data_b[21] bl[173] br[173] vss 
+ write_mux 
* No parameters

xmux_174 
+ we[6] data[21] data_b[21] bl[174] br[174] vss 
+ write_mux 
* No parameters

xmux_175 
+ we[7] data[21] data_b[21] bl[175] br[175] vss 
+ write_mux 
* No parameters

xmux_176 
+ we[0] data[22] data_b[22] bl[176] br[176] vss 
+ write_mux 
* No parameters

xmux_177 
+ we[1] data[22] data_b[22] bl[177] br[177] vss 
+ write_mux 
* No parameters

xmux_178 
+ we[2] data[22] data_b[22] bl[178] br[178] vss 
+ write_mux 
* No parameters

xmux_179 
+ we[3] data[22] data_b[22] bl[179] br[179] vss 
+ write_mux 
* No parameters

xmux_180 
+ we[4] data[22] data_b[22] bl[180] br[180] vss 
+ write_mux 
* No parameters

xmux_181 
+ we[5] data[22] data_b[22] bl[181] br[181] vss 
+ write_mux 
* No parameters

xmux_182 
+ we[6] data[22] data_b[22] bl[182] br[182] vss 
+ write_mux 
* No parameters

xmux_183 
+ we[7] data[22] data_b[22] bl[183] br[183] vss 
+ write_mux 
* No parameters

xmux_184 
+ we[0] data[23] data_b[23] bl[184] br[184] vss 
+ write_mux 
* No parameters

xmux_185 
+ we[1] data[23] data_b[23] bl[185] br[185] vss 
+ write_mux 
* No parameters

xmux_186 
+ we[2] data[23] data_b[23] bl[186] br[186] vss 
+ write_mux 
* No parameters

xmux_187 
+ we[3] data[23] data_b[23] bl[187] br[187] vss 
+ write_mux 
* No parameters

xmux_188 
+ we[4] data[23] data_b[23] bl[188] br[188] vss 
+ write_mux 
* No parameters

xmux_189 
+ we[5] data[23] data_b[23] bl[189] br[189] vss 
+ write_mux 
* No parameters

xmux_190 
+ we[6] data[23] data_b[23] bl[190] br[190] vss 
+ write_mux 
* No parameters

xmux_191 
+ we[7] data[23] data_b[23] bl[191] br[191] vss 
+ write_mux 
* No parameters

xmux_192 
+ we[0] data[24] data_b[24] bl[192] br[192] vss 
+ write_mux 
* No parameters

xmux_193 
+ we[1] data[24] data_b[24] bl[193] br[193] vss 
+ write_mux 
* No parameters

xmux_194 
+ we[2] data[24] data_b[24] bl[194] br[194] vss 
+ write_mux 
* No parameters

xmux_195 
+ we[3] data[24] data_b[24] bl[195] br[195] vss 
+ write_mux 
* No parameters

xmux_196 
+ we[4] data[24] data_b[24] bl[196] br[196] vss 
+ write_mux 
* No parameters

xmux_197 
+ we[5] data[24] data_b[24] bl[197] br[197] vss 
+ write_mux 
* No parameters

xmux_198 
+ we[6] data[24] data_b[24] bl[198] br[198] vss 
+ write_mux 
* No parameters

xmux_199 
+ we[7] data[24] data_b[24] bl[199] br[199] vss 
+ write_mux 
* No parameters

xmux_200 
+ we[0] data[25] data_b[25] bl[200] br[200] vss 
+ write_mux 
* No parameters

xmux_201 
+ we[1] data[25] data_b[25] bl[201] br[201] vss 
+ write_mux 
* No parameters

xmux_202 
+ we[2] data[25] data_b[25] bl[202] br[202] vss 
+ write_mux 
* No parameters

xmux_203 
+ we[3] data[25] data_b[25] bl[203] br[203] vss 
+ write_mux 
* No parameters

xmux_204 
+ we[4] data[25] data_b[25] bl[204] br[204] vss 
+ write_mux 
* No parameters

xmux_205 
+ we[5] data[25] data_b[25] bl[205] br[205] vss 
+ write_mux 
* No parameters

xmux_206 
+ we[6] data[25] data_b[25] bl[206] br[206] vss 
+ write_mux 
* No parameters

xmux_207 
+ we[7] data[25] data_b[25] bl[207] br[207] vss 
+ write_mux 
* No parameters

xmux_208 
+ we[0] data[26] data_b[26] bl[208] br[208] vss 
+ write_mux 
* No parameters

xmux_209 
+ we[1] data[26] data_b[26] bl[209] br[209] vss 
+ write_mux 
* No parameters

xmux_210 
+ we[2] data[26] data_b[26] bl[210] br[210] vss 
+ write_mux 
* No parameters

xmux_211 
+ we[3] data[26] data_b[26] bl[211] br[211] vss 
+ write_mux 
* No parameters

xmux_212 
+ we[4] data[26] data_b[26] bl[212] br[212] vss 
+ write_mux 
* No parameters

xmux_213 
+ we[5] data[26] data_b[26] bl[213] br[213] vss 
+ write_mux 
* No parameters

xmux_214 
+ we[6] data[26] data_b[26] bl[214] br[214] vss 
+ write_mux 
* No parameters

xmux_215 
+ we[7] data[26] data_b[26] bl[215] br[215] vss 
+ write_mux 
* No parameters

xmux_216 
+ we[0] data[27] data_b[27] bl[216] br[216] vss 
+ write_mux 
* No parameters

xmux_217 
+ we[1] data[27] data_b[27] bl[217] br[217] vss 
+ write_mux 
* No parameters

xmux_218 
+ we[2] data[27] data_b[27] bl[218] br[218] vss 
+ write_mux 
* No parameters

xmux_219 
+ we[3] data[27] data_b[27] bl[219] br[219] vss 
+ write_mux 
* No parameters

xmux_220 
+ we[4] data[27] data_b[27] bl[220] br[220] vss 
+ write_mux 
* No parameters

xmux_221 
+ we[5] data[27] data_b[27] bl[221] br[221] vss 
+ write_mux 
* No parameters

xmux_222 
+ we[6] data[27] data_b[27] bl[222] br[222] vss 
+ write_mux 
* No parameters

xmux_223 
+ we[7] data[27] data_b[27] bl[223] br[223] vss 
+ write_mux 
* No parameters

xmux_224 
+ we[0] data[28] data_b[28] bl[224] br[224] vss 
+ write_mux 
* No parameters

xmux_225 
+ we[1] data[28] data_b[28] bl[225] br[225] vss 
+ write_mux 
* No parameters

xmux_226 
+ we[2] data[28] data_b[28] bl[226] br[226] vss 
+ write_mux 
* No parameters

xmux_227 
+ we[3] data[28] data_b[28] bl[227] br[227] vss 
+ write_mux 
* No parameters

xmux_228 
+ we[4] data[28] data_b[28] bl[228] br[228] vss 
+ write_mux 
* No parameters

xmux_229 
+ we[5] data[28] data_b[28] bl[229] br[229] vss 
+ write_mux 
* No parameters

xmux_230 
+ we[6] data[28] data_b[28] bl[230] br[230] vss 
+ write_mux 
* No parameters

xmux_231 
+ we[7] data[28] data_b[28] bl[231] br[231] vss 
+ write_mux 
* No parameters

xmux_232 
+ we[0] data[29] data_b[29] bl[232] br[232] vss 
+ write_mux 
* No parameters

xmux_233 
+ we[1] data[29] data_b[29] bl[233] br[233] vss 
+ write_mux 
* No parameters

xmux_234 
+ we[2] data[29] data_b[29] bl[234] br[234] vss 
+ write_mux 
* No parameters

xmux_235 
+ we[3] data[29] data_b[29] bl[235] br[235] vss 
+ write_mux 
* No parameters

xmux_236 
+ we[4] data[29] data_b[29] bl[236] br[236] vss 
+ write_mux 
* No parameters

xmux_237 
+ we[5] data[29] data_b[29] bl[237] br[237] vss 
+ write_mux 
* No parameters

xmux_238 
+ we[6] data[29] data_b[29] bl[238] br[238] vss 
+ write_mux 
* No parameters

xmux_239 
+ we[7] data[29] data_b[29] bl[239] br[239] vss 
+ write_mux 
* No parameters

xmux_240 
+ we[0] data[30] data_b[30] bl[240] br[240] vss 
+ write_mux 
* No parameters

xmux_241 
+ we[1] data[30] data_b[30] bl[241] br[241] vss 
+ write_mux 
* No parameters

xmux_242 
+ we[2] data[30] data_b[30] bl[242] br[242] vss 
+ write_mux 
* No parameters

xmux_243 
+ we[3] data[30] data_b[30] bl[243] br[243] vss 
+ write_mux 
* No parameters

xmux_244 
+ we[4] data[30] data_b[30] bl[244] br[244] vss 
+ write_mux 
* No parameters

xmux_245 
+ we[5] data[30] data_b[30] bl[245] br[245] vss 
+ write_mux 
* No parameters

xmux_246 
+ we[6] data[30] data_b[30] bl[246] br[246] vss 
+ write_mux 
* No parameters

xmux_247 
+ we[7] data[30] data_b[30] bl[247] br[247] vss 
+ write_mux 
* No parameters

xmux_248 
+ we[0] data[31] data_b[31] bl[248] br[248] vss 
+ write_mux 
* No parameters

xmux_249 
+ we[1] data[31] data_b[31] bl[249] br[249] vss 
+ write_mux 
* No parameters

xmux_250 
+ we[2] data[31] data_b[31] bl[250] br[250] vss 
+ write_mux 
* No parameters

xmux_251 
+ we[3] data[31] data_b[31] bl[251] br[251] vss 
+ write_mux 
* No parameters

xmux_252 
+ we[4] data[31] data_b[31] bl[252] br[252] vss 
+ write_mux 
* No parameters

xmux_253 
+ we[5] data[31] data_b[31] bl[253] br[253] vss 
+ write_mux 
* No parameters

xmux_254 
+ we[6] data[31] data_b[31] bl[254] br[254] vss 
+ write_mux 
* No parameters

xmux_255 
+ we[7] data[31] data_b[31] bl[255] br[255] vss 
+ write_mux 
* No parameters

.ENDS

.SUBCKT data_dff_array 
+ vdd vss clk d[31] d[30] d[29] d[28] d[27] d[26] d[25] d[24] d[23] d[22] d[21] d[20] d[19] d[18] d[17] d[16] d[15] d[14] d[13] d[12] d[11] d[10] d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[31] q[30] q[29] q[28] q[27] q[26] q[25] q[24] q[23] q[22] q[21] q[20] q[19] q[18] q[17] q[16] q[15] q[14] q[13] q[12] q[11] q[10] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[31] q_b[30] q_b[29] q_b[28] q_b[27] q_b[26] q_b[25] q_b[24] q_b[23] q_b[22] q_b[21] q_b[20] q_b[19] q_b[18] q_b[17] q_b[16] q_b[15] q_b[14] q_b[13] q_b[12] q_b[11] q_b[10] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

xdff_10 
+ vdd vss clk d[10] q[10] q_b[10] 
+ openram_dff 
* No parameters

xdff_11 
+ vdd vss clk d[11] q[11] q_b[11] 
+ openram_dff 
* No parameters

xdff_12 
+ vdd vss clk d[12] q[12] q_b[12] 
+ openram_dff 
* No parameters

xdff_13 
+ vdd vss clk d[13] q[13] q_b[13] 
+ openram_dff 
* No parameters

xdff_14 
+ vdd vss clk d[14] q[14] q_b[14] 
+ openram_dff 
* No parameters

xdff_15 
+ vdd vss clk d[15] q[15] q_b[15] 
+ openram_dff 
* No parameters

xdff_16 
+ vdd vss clk d[16] q[16] q_b[16] 
+ openram_dff 
* No parameters

xdff_17 
+ vdd vss clk d[17] q[17] q_b[17] 
+ openram_dff 
* No parameters

xdff_18 
+ vdd vss clk d[18] q[18] q_b[18] 
+ openram_dff 
* No parameters

xdff_19 
+ vdd vss clk d[19] q[19] q_b[19] 
+ openram_dff 
* No parameters

xdff_20 
+ vdd vss clk d[20] q[20] q_b[20] 
+ openram_dff 
* No parameters

xdff_21 
+ vdd vss clk d[21] q[21] q_b[21] 
+ openram_dff 
* No parameters

xdff_22 
+ vdd vss clk d[22] q[22] q_b[22] 
+ openram_dff 
* No parameters

xdff_23 
+ vdd vss clk d[23] q[23] q_b[23] 
+ openram_dff 
* No parameters

xdff_24 
+ vdd vss clk d[24] q[24] q_b[24] 
+ openram_dff 
* No parameters

xdff_25 
+ vdd vss clk d[25] q[25] q_b[25] 
+ openram_dff 
* No parameters

xdff_26 
+ vdd vss clk d[26] q[26] q_b[26] 
+ openram_dff 
* No parameters

xdff_27 
+ vdd vss clk d[27] q[27] q_b[27] 
+ openram_dff 
* No parameters

xdff_28 
+ vdd vss clk d[28] q[28] q_b[28] 
+ openram_dff 
* No parameters

xdff_29 
+ vdd vss clk d[29] q[29] q_b[29] 
+ openram_dff 
* No parameters

xdff_30 
+ vdd vss clk d[30] q[30] q_b[30] 
+ openram_dff 
* No parameters

xdff_31 
+ vdd vss clk d[31] q[31] q_b[31] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT addr_dff_array 
+ vdd vss clk d[4] d[3] d[2] d[1] d[0] q[4] q[3] q[2] q[1] q[0] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT col_data_inv 
+ din din_b vdd vss 

xMP0 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.6' l='0.15' 

xMN0 
+ din_b din vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.4' l='0.15' 

.ENDS

.SUBCKT col_inv_array 
+ din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] din_b[31] din_b[30] din_b[29] din_b[28] din_b[27] din_b[26] din_b[25] din_b[24] din_b[23] din_b[22] din_b[21] din_b[20] din_b[19] din_b[18] din_b[17] din_b[16] din_b[15] din_b[14] din_b[13] din_b[12] din_b[11] din_b[10] din_b[9] din_b[8] din_b[7] din_b[6] din_b[5] din_b[4] din_b[3] din_b[2] din_b[1] din_b[0] vdd vss 

xinv_0 
+ din[0] din_b[0] vdd vss 
+ col_data_inv 
* No parameters

xinv_1 
+ din[1] din_b[1] vdd vss 
+ col_data_inv 
* No parameters

xinv_2 
+ din[2] din_b[2] vdd vss 
+ col_data_inv 
* No parameters

xinv_3 
+ din[3] din_b[3] vdd vss 
+ col_data_inv 
* No parameters

xinv_4 
+ din[4] din_b[4] vdd vss 
+ col_data_inv 
* No parameters

xinv_5 
+ din[5] din_b[5] vdd vss 
+ col_data_inv 
* No parameters

xinv_6 
+ din[6] din_b[6] vdd vss 
+ col_data_inv 
* No parameters

xinv_7 
+ din[7] din_b[7] vdd vss 
+ col_data_inv 
* No parameters

xinv_8 
+ din[8] din_b[8] vdd vss 
+ col_data_inv 
* No parameters

xinv_9 
+ din[9] din_b[9] vdd vss 
+ col_data_inv 
* No parameters

xinv_10 
+ din[10] din_b[10] vdd vss 
+ col_data_inv 
* No parameters

xinv_11 
+ din[11] din_b[11] vdd vss 
+ col_data_inv 
* No parameters

xinv_12 
+ din[12] din_b[12] vdd vss 
+ col_data_inv 
* No parameters

xinv_13 
+ din[13] din_b[13] vdd vss 
+ col_data_inv 
* No parameters

xinv_14 
+ din[14] din_b[14] vdd vss 
+ col_data_inv 
* No parameters

xinv_15 
+ din[15] din_b[15] vdd vss 
+ col_data_inv 
* No parameters

xinv_16 
+ din[16] din_b[16] vdd vss 
+ col_data_inv 
* No parameters

xinv_17 
+ din[17] din_b[17] vdd vss 
+ col_data_inv 
* No parameters

xinv_18 
+ din[18] din_b[18] vdd vss 
+ col_data_inv 
* No parameters

xinv_19 
+ din[19] din_b[19] vdd vss 
+ col_data_inv 
* No parameters

xinv_20 
+ din[20] din_b[20] vdd vss 
+ col_data_inv 
* No parameters

xinv_21 
+ din[21] din_b[21] vdd vss 
+ col_data_inv 
* No parameters

xinv_22 
+ din[22] din_b[22] vdd vss 
+ col_data_inv 
* No parameters

xinv_23 
+ din[23] din_b[23] vdd vss 
+ col_data_inv 
* No parameters

xinv_24 
+ din[24] din_b[24] vdd vss 
+ col_data_inv 
* No parameters

xinv_25 
+ din[25] din_b[25] vdd vss 
+ col_data_inv 
* No parameters

xinv_26 
+ din[26] din_b[26] vdd vss 
+ col_data_inv 
* No parameters

xinv_27 
+ din[27] din_b[27] vdd vss 
+ col_data_inv 
* No parameters

xinv_28 
+ din[28] din_b[28] vdd vss 
+ col_data_inv 
* No parameters

xinv_29 
+ din[29] din_b[29] vdd vss 
+ col_data_inv 
* No parameters

xinv_30 
+ din[30] din_b[30] vdd vss 
+ col_data_inv 
* No parameters

xinv_31 
+ din[31] din_b[31] vdd vss 
+ col_data_inv 
* No parameters

.ENDS

.SUBCKT sense_amp_array 
+ vdd vss clk bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] 

xsense_amp_0 
+ clk br[0] bl[0] data_b[0] data[0] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_1 
+ clk br[1] bl[1] data_b[1] data[1] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_2 
+ clk br[2] bl[2] data_b[2] data[2] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_3 
+ clk br[3] bl[3] data_b[3] data[3] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_4 
+ clk br[4] bl[4] data_b[4] data[4] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_5 
+ clk br[5] bl[5] data_b[5] data[5] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_6 
+ clk br[6] bl[6] data_b[6] data[6] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_7 
+ clk br[7] bl[7] data_b[7] data[7] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_8 
+ clk br[8] bl[8] data_b[8] data[8] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_9 
+ clk br[9] bl[9] data_b[9] data[9] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_10 
+ clk br[10] bl[10] data_b[10] data[10] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_11 
+ clk br[11] bl[11] data_b[11] data[11] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_12 
+ clk br[12] bl[12] data_b[12] data[12] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_13 
+ clk br[13] bl[13] data_b[13] data[13] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_14 
+ clk br[14] bl[14] data_b[14] data[14] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_15 
+ clk br[15] bl[15] data_b[15] data[15] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_16 
+ clk br[16] bl[16] data_b[16] data[16] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_17 
+ clk br[17] bl[17] data_b[17] data[17] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_18 
+ clk br[18] bl[18] data_b[18] data[18] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_19 
+ clk br[19] bl[19] data_b[19] data[19] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_20 
+ clk br[20] bl[20] data_b[20] data[20] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_21 
+ clk br[21] bl[21] data_b[21] data[21] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_22 
+ clk br[22] bl[22] data_b[22] data[22] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_23 
+ clk br[23] bl[23] data_b[23] data[23] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_24 
+ clk br[24] bl[24] data_b[24] data[24] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_25 
+ clk br[25] bl[25] data_b[25] data[25] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_26 
+ clk br[26] bl[26] data_b[26] data[26] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_27 
+ clk br[27] bl[27] data_b[27] data[27] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_28 
+ clk br[28] bl[28] data_b[28] data[28] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_29 
+ clk br[29] bl[29] data_b[29] data[29] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_30 
+ clk br[30] bl[30] data_b[30] data[30] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_31 
+ clk br[31] bl[31] data_b[31] data[31] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

.ENDS

.SUBCKT dout_buf 
+ din1 din2 dout1 dout2 vdd vss 

xMP11 
+ x1 din1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN11 
+ x1 din1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP21 
+ dout1 x1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN21 
+ dout1 x1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMP12 
+ x2 din2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN12 
+ x2 din2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP22 
+ dout2 x2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN22 
+ dout2 x2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dout_buf_array 
+ din1[31] din1[30] din1[29] din1[28] din1[27] din1[26] din1[25] din1[24] din1[23] din1[22] din1[21] din1[20] din1[19] din1[18] din1[17] din1[16] din1[15] din1[14] din1[13] din1[12] din1[11] din1[10] din1[9] din1[8] din1[7] din1[6] din1[5] din1[4] din1[3] din1[2] din1[1] din1[0] din2[31] din2[30] din2[29] din2[28] din2[27] din2[26] din2[25] din2[24] din2[23] din2[22] din2[21] din2[20] din2[19] din2[18] din2[17] din2[16] din2[15] din2[14] din2[13] din2[12] din2[11] din2[10] din2[9] din2[8] din2[7] din2[6] din2[5] din2[4] din2[3] din2[2] din2[1] din2[0] dout1[31] dout1[30] dout1[29] dout1[28] dout1[27] dout1[26] dout1[25] dout1[24] dout1[23] dout1[22] dout1[21] dout1[20] dout1[19] dout1[18] dout1[17] dout1[16] dout1[15] dout1[14] dout1[13] dout1[12] dout1[11] dout1[10] dout1[9] dout1[8] dout1[7] dout1[6] dout1[5] dout1[4] dout1[3] dout1[2] dout1[1] dout1[0] dout2[31] dout2[30] dout2[29] dout2[28] dout2[27] dout2[26] dout2[25] dout2[24] dout2[23] dout2[22] dout2[21] dout2[20] dout2[19] dout2[18] dout2[17] dout2[16] dout2[15] dout2[14] dout2[13] dout2[12] dout2[11] dout2[10] dout2[9] dout2[8] dout2[7] dout2[6] dout2[5] dout2[4] dout2[3] dout2[2] dout2[1] dout2[0] vdd vss 

xbuf_0 
+ din1[0] din2[0] dout1[0] dout2[0] vdd vss 
+ dout_buf 
* No parameters

xbuf_1 
+ din1[1] din2[1] dout1[1] dout2[1] vdd vss 
+ dout_buf 
* No parameters

xbuf_2 
+ din1[2] din2[2] dout1[2] dout2[2] vdd vss 
+ dout_buf 
* No parameters

xbuf_3 
+ din1[3] din2[3] dout1[3] dout2[3] vdd vss 
+ dout_buf 
* No parameters

xbuf_4 
+ din1[4] din2[4] dout1[4] dout2[4] vdd vss 
+ dout_buf 
* No parameters

xbuf_5 
+ din1[5] din2[5] dout1[5] dout2[5] vdd vss 
+ dout_buf 
* No parameters

xbuf_6 
+ din1[6] din2[6] dout1[6] dout2[6] vdd vss 
+ dout_buf 
* No parameters

xbuf_7 
+ din1[7] din2[7] dout1[7] dout2[7] vdd vss 
+ dout_buf 
* No parameters

xbuf_8 
+ din1[8] din2[8] dout1[8] dout2[8] vdd vss 
+ dout_buf 
* No parameters

xbuf_9 
+ din1[9] din2[9] dout1[9] dout2[9] vdd vss 
+ dout_buf 
* No parameters

xbuf_10 
+ din1[10] din2[10] dout1[10] dout2[10] vdd vss 
+ dout_buf 
* No parameters

xbuf_11 
+ din1[11] din2[11] dout1[11] dout2[11] vdd vss 
+ dout_buf 
* No parameters

xbuf_12 
+ din1[12] din2[12] dout1[12] dout2[12] vdd vss 
+ dout_buf 
* No parameters

xbuf_13 
+ din1[13] din2[13] dout1[13] dout2[13] vdd vss 
+ dout_buf 
* No parameters

xbuf_14 
+ din1[14] din2[14] dout1[14] dout2[14] vdd vss 
+ dout_buf 
* No parameters

xbuf_15 
+ din1[15] din2[15] dout1[15] dout2[15] vdd vss 
+ dout_buf 
* No parameters

xbuf_16 
+ din1[16] din2[16] dout1[16] dout2[16] vdd vss 
+ dout_buf 
* No parameters

xbuf_17 
+ din1[17] din2[17] dout1[17] dout2[17] vdd vss 
+ dout_buf 
* No parameters

xbuf_18 
+ din1[18] din2[18] dout1[18] dout2[18] vdd vss 
+ dout_buf 
* No parameters

xbuf_19 
+ din1[19] din2[19] dout1[19] dout2[19] vdd vss 
+ dout_buf 
* No parameters

xbuf_20 
+ din1[20] din2[20] dout1[20] dout2[20] vdd vss 
+ dout_buf 
* No parameters

xbuf_21 
+ din1[21] din2[21] dout1[21] dout2[21] vdd vss 
+ dout_buf 
* No parameters

xbuf_22 
+ din1[22] din2[22] dout1[22] dout2[22] vdd vss 
+ dout_buf 
* No parameters

xbuf_23 
+ din1[23] din2[23] dout1[23] dout2[23] vdd vss 
+ dout_buf 
* No parameters

xbuf_24 
+ din1[24] din2[24] dout1[24] dout2[24] vdd vss 
+ dout_buf 
* No parameters

xbuf_25 
+ din1[25] din2[25] dout1[25] dout2[25] vdd vss 
+ dout_buf 
* No parameters

xbuf_26 
+ din1[26] din2[26] dout1[26] dout2[26] vdd vss 
+ dout_buf 
* No parameters

xbuf_27 
+ din1[27] din2[27] dout1[27] dout2[27] vdd vss 
+ dout_buf 
* No parameters

xbuf_28 
+ din1[28] din2[28] dout1[28] dout2[28] vdd vss 
+ dout_buf 
* No parameters

xbuf_29 
+ din1[29] din2[29] dout1[29] dout2[29] vdd vss 
+ dout_buf 
* No parameters

xbuf_30 
+ din1[30] din2[30] dout1[30] dout2[30] vdd vss 
+ dout_buf 
* No parameters

xbuf_31 
+ din1[31] din2[31] dout1[31] dout2[31] vdd vss 
+ dout_buf 
* No parameters

.ENDS

.SUBCKT we_control_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='8.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='12.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ we_control_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ we_control_and2_inv 
* No parameters

.ENDS

.SUBCKT we_control 
+ wr_en sel[7] sel[6] sel[5] sel[4] sel[3] sel[2] sel[1] sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 

xand2_0 
+ sel[0] wr_en write_driver_en[0] vdd vss 
+ we_control_and2 
* No parameters

xand2_1 
+ sel[1] wr_en write_driver_en[1] vdd vss 
+ we_control_and2 
* No parameters

xand2_2 
+ sel[2] wr_en write_driver_en[2] vdd vss 
+ we_control_and2 
* No parameters

xand2_3 
+ sel[3] wr_en write_driver_en[3] vdd vss 
+ we_control_and2 
* No parameters

xand2_4 
+ sel[4] wr_en write_driver_en[4] vdd vss 
+ we_control_and2 
* No parameters

xand2_5 
+ sel[5] wr_en write_driver_en[5] vdd vss 
+ we_control_and2 
* No parameters

xand2_6 
+ sel[6] wr_en write_driver_en[6] vdd vss 
+ we_control_and2 
* No parameters

xand2_7 
+ sel[7] wr_en write_driver_en[7] vdd vss 
+ we_control_and2 
* No parameters

.ENDS

.SUBCKT control_logic_delay_chain 
+ din dout vdd vss 

xinv_0 
+ din int[0] vdd vss 
+ control_logic_inv 
* No parameters

xinv_1 
+ int[0] int[1] vdd vss 
+ control_logic_inv 
* No parameters

xinv_2 
+ int[1] int[2] vdd vss 
+ control_logic_inv 
* No parameters

xinv_3 
+ int[2] int[3] vdd vss 
+ control_logic_inv 
* No parameters

xinv_4 
+ int[3] int[4] vdd vss 
+ control_logic_inv 
* No parameters

xinv_5 
+ int[4] int[5] vdd vss 
+ control_logic_inv 
* No parameters

xinv_6 
+ int[5] int[6] vdd vss 
+ control_logic_inv 
* No parameters

xinv_7 
+ int[6] int[7] vdd vss 
+ control_logic_inv 
* No parameters

xinv_8 
+ int[7] int[8] vdd vss 
+ control_logic_inv 
* No parameters

xinv_9 
+ int[8] int[9] vdd vss 
+ control_logic_inv 
* No parameters

xinv_10 
+ int[9] int[10] vdd vss 
+ control_logic_inv 
* No parameters

xinv_11 
+ int[10] int[11] vdd vss 
+ control_logic_inv 
* No parameters

xinv_12 
+ int[11] int[12] vdd vss 
+ control_logic_inv 
* No parameters

xinv_13 
+ int[12] int[13] vdd vss 
+ control_logic_inv 
* No parameters

xinv_14 
+ int[13] int[14] vdd vss 
+ control_logic_inv 
* No parameters

xinv_15 
+ int[14] int[15] vdd vss 
+ control_logic_inv 
* No parameters

xinv_16 
+ int[15] int[16] vdd vss 
+ control_logic_inv 
* No parameters

xinv_17 
+ int[16] int[17] vdd vss 
+ control_logic_inv 
* No parameters

xinv_18 
+ int[17] int[18] vdd vss 
+ control_logic_inv 
* No parameters

xinv_19 
+ int[18] int[19] vdd vss 
+ control_logic_inv 
* No parameters

xinv_20 
+ int[19] int[20] vdd vss 
+ control_logic_inv 
* No parameters

xinv_21 
+ int[20] int[21] vdd vss 
+ control_logic_inv 
* No parameters

xinv_22 
+ int[21] int[22] vdd vss 
+ control_logic_inv 
* No parameters

xinv_23 
+ int[22] int[23] vdd vss 
+ control_logic_inv 
* No parameters

xinv_24 
+ int[23] int[24] vdd vss 
+ control_logic_inv 
* No parameters

xinv_25 
+ int[24] int[25] vdd vss 
+ control_logic_inv 
* No parameters

xinv_26 
+ int[25] int[26] vdd vss 
+ control_logic_inv 
* No parameters

xinv_27 
+ int[26] int[27] vdd vss 
+ control_logic_inv 
* No parameters

xinv_28 
+ int[27] int[28] vdd vss 
+ control_logic_inv 
* No parameters

xinv_29 
+ int[28] int[29] vdd vss 
+ control_logic_inv 
* No parameters

xinv_30 
+ int[29] int[30] vdd vss 
+ control_logic_inv 
* No parameters

xinv_31 
+ int[30] int[31] vdd vss 
+ control_logic_inv 
* No parameters

xinv_32 
+ int[31] int[32] vdd vss 
+ control_logic_inv 
* No parameters

xinv_33 
+ int[32] int[33] vdd vss 
+ control_logic_inv 
* No parameters

xinv_34 
+ int[33] int[34] vdd vss 
+ control_logic_inv 
* No parameters

xinv_35 
+ int[34] int[35] vdd vss 
+ control_logic_inv 
* No parameters

xinv_36 
+ int[35] int[36] vdd vss 
+ control_logic_inv 
* No parameters

xinv_37 
+ int[36] int[37] vdd vss 
+ control_logic_inv 
* No parameters

xinv_38 
+ int[37] int[38] vdd vss 
+ control_logic_inv 
* No parameters

xinv_39 
+ int[38] int[39] vdd vss 
+ control_logic_inv 
* No parameters

xinv_40 
+ int[39] int[40] vdd vss 
+ control_logic_inv 
* No parameters

xinv_41 
+ int[40] int[41] vdd vss 
+ control_logic_inv 
* No parameters

xinv_42 
+ int[41] int[42] vdd vss 
+ control_logic_inv 
* No parameters

xinv_43 
+ int[42] int[43] vdd vss 
+ control_logic_inv 
* No parameters

xinv_44 
+ int[43] dout vdd vss 
+ control_logic_inv 
* No parameters

.ENDS

.SUBCKT sramgen_sram_32x32m8w32_replica_v1 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] we addr[4] addr[3] addr[2] addr[1] addr[0] 

xdin_dffs 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] dff_din_b[31] dff_din_b[30] dff_din_b[29] dff_din_b[28] dff_din_b[27] dff_din_b[26] dff_din_b[25] dff_din_b[24] dff_din_b[23] dff_din_b[22] dff_din_b[21] dff_din_b[20] dff_din_b[19] dff_din_b[18] dff_din_b[17] dff_din_b[16] dff_din_b[15] dff_din_b[14] dff_din_b[13] dff_din_b[12] dff_din_b[11] dff_din_b[10] dff_din_b[9] dff_din_b[8] dff_din_b[7] dff_din_b[6] dff_din_b[5] dff_din_b[4] dff_din_b[3] dff_din_b[2] dff_din_b[1] dff_din_b[0] 
+ data_dff_array 
* No parameters

xaddr_dffs 
+ vdd vss clk addr[4] addr[3] addr[2] addr[1] addr[0] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] 
+ addr_dff_array 
* No parameters

xwe_dff 
+ vdd vss clk we bank_we bank_we_b 
+ openram_dff 
* No parameters

xdecoder 
+ vdd vss bank_addr[4] bank_addr[3] bank_addr_b[4] bank_addr_b[3] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_data_b[3] wl_data_b[2] wl_data_b[1] wl_data_b[0] 
+ hierarchical_decoder 
* No parameters

xwl_driver_array 
+ vdd vss wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_en wl[3] wl[2] wl[1] wl[0] 
+ wordline_driver_array 
* No parameters

xbitcells 
+ vdd vss bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[3] wl[2] wl[1] wl[0] vss vdd rbl rbr 
+ bitcell_array 
* No parameters

xprecharge_array 
+ vdd pc_b rbl bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0]  rbr br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0]  
+ precharge_array 
* No parameters

xwrite_mux_array 
+ write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 
+ write_mux_array 
* No parameters

xread_mux_array 
+ col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] vdd 
+ read_mux_array 
* No parameters

xcol_inv_array 
+ bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] vdd vss 
+ col_inv_array 
* No parameters

xsense_amp_array 
+ vdd vss sense_amp_en bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] 
+ sense_amp_array 
* No parameters

xdout_buf_array 
+ sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] dout_b[31] dout_b[30] dout_b[29] dout_b[28] dout_b[27] dout_b[26] dout_b[25] dout_b[24] dout_b[23] dout_b[22] dout_b[21] dout_b[20] dout_b[19] dout_b[18] dout_b[17] dout_b[16] dout_b[15] dout_b[14] dout_b[13] dout_b[12] dout_b[11] dout_b[10] dout_b[9] dout_b[8] dout_b[7] dout_b[6] dout_b[5] dout_b[4] dout_b[3] dout_b[2] dout_b[1] dout_b[0] vdd vss 
+ dout_buf_array 
* No parameters

xcontrol_logic 
+ clk bank_we rbl pc_b wl_en wr_en sense_amp_en vdd vss 
+ sramgen_control_replica_v1 
* No parameters

xcolumn_decoder 
+ vdd vss bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] 
+ column_decoder 
* No parameters

xwe_control 
+ wr_en col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 
+ we_control 
* No parameters

.ENDS

